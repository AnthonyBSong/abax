module vvadd_mem(
  input wire clk,
  input wire rst,
  input wire out_rdy,
  input wire v0__read_req_rdy,
  input wire [31:0] v0__read_resp,
  input wire v0__read_resp_vld,
  input wire v0__write_completion_vld,
  input wire v0__write_req_rdy,
  input wire [31:0] v0_in,
  input wire v0_in_vld,
  input wire v1__read_req_rdy,
  input wire [31:0] v1__read_resp,
  input wire v1__read_resp_vld,
  input wire v1__write_completion_vld,
  input wire v1__write_req_rdy,
  input wire [31:0] v1_in,
  input wire v1_in_vld,
  input wire [31:0] c_rd_data,
  output wire [31:0] out,
  output wire out_vld,
  output wire [3:0] v0__read_req,
  output wire v0__read_req_vld,
  output wire v0__read_resp_rdy,
  output wire v0__write_completion_rdy,
  output wire [35:0] v0__write_req,
  output wire v0__write_req_vld,
  output wire v0_in_rdy,
  output wire [3:0] v1__read_req,
  output wire v1__read_req_vld,
  output wire v1__read_resp_rdy,
  output wire v1__write_completion_rdy,
  output wire [35:0] v1__write_req,
  output wire v1__write_req_vld,
  output wire v1_in_rdy,
  output wire [3:0] c_rd_addr,
  output wire c_rd_en,
  output wire [3:0] c_wr_addr,
  output wire [31:0] c_wr_data,
  output wire c_wr_en
);
  wire [31:0] literal_11058 = 32'h0000_0000;
  wire [31:0] literal_11062 = 32'h0000_0000;
  wire [31:0] literal_11126 = 32'h0000_0000;
  reg ____for_1__last_iter_broke;
  reg [1:0] __this_1;
  reg [4:0] ____for_1_i;
  reg [31:0] __this_0;
  reg ____fsm_vvadd_impl_state_2;
  reg [4:0] ____fsm_vvadd_impl_state_0;
  reg ____fsm_vvadd_impl_state_4;
  reg ____fsm_vvadd_impl_exited_last_activation;
  reg [4:0] p0_____fsm_vvadd_impl_state_0__1;
  reg p0___fsm_vvadd_impl_in_state_0;
  reg p0_continuation_9_ctx_4__relative_c_output;
  reg p0___for_1_loop_contents_condition;
  reg p0_nor_10933;
  reg p0_and_10968;
  reg p0_and_10971;
  reg p0_nand_10999;
  reg p0_and_10903;
  reg p0_and_10904;
  reg p0_and_10905;
  reg p0_and_10906;
  reg p1___for_1_loop_contents_condition;
  reg p1_and_11120;
  reg p1_and_11090;
  reg p1_and_11089;
  reg p1_and_11076;
  reg p1_and_11087;
  reg p1_and_11072;
  reg p1_and_11070;
  reg p1_and_11054;
  reg p1_and_11084;
  reg p1_and_11083;
  reg p1_and_11082;
  reg p1_and_11075;
  reg p1_and_11081;
  reg p1_and_11071;
  reg p1_and_11069;
  reg p1_and_11053;
  reg p1_or_11123;
  reg p1_nand_10999;
  reg p1_nand_11132;
  reg p1_nand_11133;
  reg p1_nand_11134;
  reg p1_nand_11135;
  reg p1_nand_11136;
  reg p1_nand_11137;
  reg p1_nand_11138;
  reg p1_nand_11139;
  reg p1_nand_11140;
  reg p1_nand_11141;
  reg p1_nand_11142;
  reg p1_nand_11143;
  reg p1_nand_11144;
  reg p1_nand_11145;
  reg p1_nand_11146;
  reg p1_nand_11147;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg p4_valid;
  reg __v0__read_req_has_been_sent_reg;
  reg __v1__read_req_has_been_sent_reg;
  reg __c__read_req_has_been_sent_reg;
  reg __v0__write_req_has_been_sent_reg;
  reg __v1__write_req_has_been_sent_reg;
  reg __c__write_req_has_been_sent_reg;
  reg __out_has_been_sent_reg;
  reg __c_rd_en__1_delay_reg;
  reg [31:0] __c_ram_zero_latency0_skid_reg;
  reg __c_ram_zero_latency0_valid_skid_reg;
  wire __fsm_vvadd_impl_default_next_state;
  wire [4:0] and_10856;
  wire [4:0] __fsm_vvadd_impl_state_0_index;
  wire __fsm_vvadd_impl_in_state_0;
  wire continuation_1_ctx_3__full_condi_output__1;
  wire eq_10859;
  wire [5:0] add_10862;
  wire [1:0] unexpand_for_this_next_1_case_1_case_1_case_1;
  wire [1:0] unexpand_for_this_next_1_case_1_case_0_case_0_case_1;
  wire nor_10876;
  wire [1:0] sel_10864;
  wire [1:0] unexpand_for_this_next_1_case_1_case_1_case_0;
  wire __for_1_do_break_from_func;
  wire v0_in_recv_valid;
  wire continuation_9_ctx_4__relative_c_output;
  wire [4:0] __fsm_vvadd_impl_state_17_index;
  wire __for_1_not_exit_state_condition;
  wire v0_read_pred;
  wire [31:0] add_10882;
  wire __fsm_vvadd_impl_in_state_17;
  wire __fsm_vvadd_impl_go_to_next_state_in_state;
  wire nand_10891;
  wire continuation_4_ctx_3__full_condi_output__2;
  wire continuation_4_ctx_3__full_condi_output;
  wire [31:0] sel_10901;
  wire [4:0] __fsm_vvadd_impl_state_16_index;
  wire and_10936;
  wire nor_10907;
  wire eq_10909;
  wire __fsm_vvadd_impl_in_state_16;
  wire v1_in_recv_valid;
  wire [4:0] __fsm_vvadd_impl_state_15_index;
  wire [4:0] __fsm_vvadd_impl_state_7_index;
  wire and_10915;
  wire and_10917;
  wire __for_1_loop_contents_condition;
  wire nor_10933;
  wire and_10968;
  wire and_10971;
  wire [4:0] __fsm_vvadd_impl_state_14_index;
  wire [4:0] __fsm_vvadd_impl_state_6_index;
  wire [4:0] __fsm_vvadd_impl_state_13_index;
  wire [4:0] __fsm_vvadd_impl_state_5_index;
  wire __fsm_vvadd_impl_in_state_15;
  wire __fsm_vvadd_impl_in_state_7;
  wire [4:0] __fsm_vvadd_impl_state_11_index;
  wire [4:0] __fsm_vvadd_impl_state_3_index;
  wire and_10923;
  wire and_10924;
  wire and_10925;
  wire and_10926;
  wire and_10927;
  wire nor_10928;
  wire __fsm_vvadd_impl_returns_this_activation_vars;
  wire and_10930;
  wire and_10931;
  wire p1_all_active_inputs_valid;
  wire p1_all_active_outputs_ready;
  wire c__read_req_not_pred;
  wire c_ram_zero_latency0_from_skid_rdy;
  wire v0__write_req_not_pred;
  wire v1__write_req_not_pred;
  wire [4:0] __fsm_vvadd_impl_state_one;
  wire [4:0] __fsm_vvadd_impl_state_2_index;
  wire [4:0] __fsm_vvadd_impl_state_4_index;
  wire [4:0] __fsm_vvadd_impl_state_8_index;
  wire [4:0] __fsm_vvadd_impl_state_9_index;
  wire [4:0] __fsm_vvadd_impl_state_10_index;
  wire [4:0] __fsm_vvadd_impl_state_12_index;
  wire __fsm_vvadd_impl_in_state_14;
  wire __fsm_vvadd_impl_in_state_6;
  wire __fsm_vvadd_impl_in_state_13;
  wire __fsm_vvadd_impl_in_state_5;
  wire and_11053;
  wire and_11054;
  wire __fsm_vvadd_impl_in_state_11;
  wire __fsm_vvadd_impl_in_state_3;
  wire [4:0] __this_0__next_value_predicates;
  wire [1:0] ____fsm_vvadd_impl_state_0__next_value_predicates;
  wire [3:0] __this_1__next_value_predicates;
  wire p1_stage_done;
  wire p1_not_valid;
  wire __fsm_vvadd_impl_in_state_1;
  wire __fsm_vvadd_impl_in_state_2;
  wire __fsm_vvadd_impl_in_state_4;
  wire __fsm_vvadd_impl_in_state_8;
  wire __fsm_vvadd_impl_in_state_9;
  wire __fsm_vvadd_impl_in_state_10;
  wire __fsm_vvadd_impl_in_state_12;
  wire and_11069;
  wire and_11070;
  wire and_11071;
  wire and_11072;
  wire or_11074;
  wire and_11075;
  wire and_11076;
  wire [31:0] v0__read_resp_select;
  wire [31:0] v1__read_resp_select;
  wire [5:0] one_hot_10947;
  wire [2:0] one_hot_10948;
  wire [4:0] one_hot_10949;
  wire p0_enable;
  wire p0_all_active_outputs_ready;
  wire and_11120;
  wire and_11090;
  wire and_11089;
  wire and_11087;
  wire and_11084;
  wire and_11083;
  wire and_11082;
  wire and_11081;
  wire or_11085;
  wire or_11086;
  wire or_11088;
  wire [31:0] v0_read_response;
  wire [31:0] v1_read_response;
  wire [31:0] c_ram_zero_latency0_select;
  wire p0_data_enable;
  wire __v0__read_req_vld_buf;
  wire __v0__read_req_not_has_been_sent;
  wire __v1__read_req_not_has_been_sent;
  wire __c__read_req_vld_buf;
  wire __c__read_req_not_has_been_sent;
  wire __v0__write_req_vld_buf;
  wire __v0__write_req_not_has_been_sent;
  wire __v1__write_req_vld_buf;
  wire __v1__write_req_not_has_been_sent;
  wire or_11123;
  wire __out_vld_buf;
  wire __out_not_has_been_sent;
  wire and_11437;
  wire [3:0] v0_write_addr;
  wire [31:0] c_write_value__16;
  wire and_11395;
  wire and_11396;
  wire and_11397;
  wire and_11398;
  wire and_11399;
  wire and_11406;
  wire and_11407;
  wire and_11418;
  wire and_11420;
  wire __v0__read_req_valid_and_not_has_been_sent;
  wire __v1__read_req_valid_and_not_has_been_sent;
  wire c_rd_en__1;
  wire __v0__write_req_valid_and_not_has_been_sent;
  wire __v1__write_req_valid_and_not_has_been_sent;
  wire __c__write_req_vld_buf;
  wire __c__write_req_not_has_been_sent;
  wire __out_valid_and_not_has_been_sent;
  wire c_ram_zero_latency0_to_is_not_rdy;
  wire [3:0] c_read_addr;
  wire [31:0] c__read_resp_select;
  wire [3:0] v0_read_addr;
  wire [31:0] v0_in_select;
  wire [3:0] v1_write_addr;
  wire [31:0] v1_in_select;
  wire __this_0__at_most_one_next_value;
  wire ____fsm_vvadd_impl_state_0__at_most_one_next_value;
  wire __this_1__at_most_one_next_value;
  wire [4:0] concat_11401;
  wire [31:0] ctx_3__x_literal__1;
  wire [31:0] add_10992;
  wire [1:0] concat_11409;
  wire [4:0] __fsm_vvadd_impl_state_plus_one;
  wire [3:0] concat_11423;
  wire [1:0] unexpand_for_this_next_1_case_1_case_0_case_1;
  wire __for_1_guarded_update_state_elements;
  wire __v0__read_req_valid_and_all_active_outputs_ready;
  wire __v0__read_req_valid_and_ready_txfr;
  wire __v1__read_req_valid_and_ready_txfr;
  wire __c__read_req_valid_and_all_active_outputs_ready;
  wire __c__read_req_valid_and_ready_txfr;
  wire __v0__write_req_valid_and_all_active_outputs_ready;
  wire __v0__write_req_valid_and_ready_txfr;
  wire __v1__write_req_valid_and_all_active_outputs_ready;
  wire __v1__write_req_valid_and_ready_txfr;
  wire __c__write_req_valid_and_all_active_outputs_ready;
  wire c_wr_en__1;
  wire __out_valid_and_all_active_outputs_ready;
  wire __out_valid_and_ready_txfr;
  wire c_ram_zero_latency0_skid_data_load_en;
  wire c_ram_zero_latency0_skid_valid_set_zero;
  wire [3:0] tuple_10932;
  wire [35:0] tuple_11122;
  wire [31:0] c_read_response;
  wire [3:0] tuple_10872;
  wire and_11439;
  wire or_11572;
  wire or_11574;
  wire or_11576;
  wire p4_enable;
  wire p3_enable;
  wire p2_enable;
  wire p1_enable;
  wire nand_11132;
  wire nand_11133;
  wire nand_11134;
  wire nand_11135;
  wire nand_11136;
  wire nand_11137;
  wire nand_11138;
  wire nand_11139;
  wire nand_11140;
  wire nand_11141;
  wire nand_11142;
  wire nand_11143;
  wire nand_11144;
  wire nand_11145;
  wire nand_11146;
  wire nand_11147;
  wire nand_10999;
  wire and_10903;
  wire and_10904;
  wire and_10905;
  wire and_10906;
  wire [31:0] one_hot_sel_11402;
  wire or_11403;
  wire [4:0] one_hot_sel_11410;
  wire or_11411;
  wire sel_10989;
  wire sel_10990;
  wire and_11415;
  wire [1:0] one_hot_sel_11424;
  wire or_11425;
  wire [4:0] unexpand_for___for_1_i_next__1_case_1;
  wire and_11427;
  wire __v0__read_req_not_stage_load;
  wire __v0__read_req_has_been_sent_reg_load_en;
  wire __v1__read_req_has_been_sent_reg_load_en;
  wire __c__read_req_not_stage_load;
  wire __c__read_req_has_been_sent_reg_load_en;
  wire __v0__write_req_not_stage_load;
  wire __v0__write_req_has_been_sent_reg_load_en;
  wire __v1__write_req_not_stage_load;
  wire __v1__write_req_has_been_sent_reg_load_en;
  wire __c__write_req_not_stage_load;
  wire __c__write_req_has_been_sent_reg_load_en;
  wire __out_not_stage_load;
  wire __out_has_been_sent_reg_load_en;
  wire c_ram_zero_latency0_skid_valid_load_en;
  assign __fsm_vvadd_impl_default_next_state = 1'h0;
  assign and_10856 = {5{~____for_1__last_iter_broke}} & ____for_1_i;
  assign __fsm_vvadd_impl_state_0_index = 5'h00;
  assign __fsm_vvadd_impl_in_state_0 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_0_index;
  assign continuation_1_ctx_3__full_condi_output__1 = ~(__this_1[0] | __this_1[1]);
  assign eq_10859 = __this_0 == 32'h0000_000f;
  assign add_10862 = {__fsm_vvadd_impl_default_next_state, and_10856} + 6'h01;
  assign unexpand_for_this_next_1_case_1_case_1_case_1 = 2'h1;
  assign unexpand_for_this_next_1_case_1_case_0_case_0_case_1 = 2'h0;
  assign nor_10876 = ~(__this_1[0] | __this_1[1] | ~__fsm_vvadd_impl_in_state_0);
  assign sel_10864 = ~(continuation_1_ctx_3__full_condi_output__1 & ____fsm_vvadd_impl_state_2 & eq_10859) ? __this_1 : unexpand_for_this_next_1_case_1_case_1_case_1;
  assign unexpand_for_this_next_1_case_1_case_1_case_0 = 2'h2;
  assign __for_1_do_break_from_func = add_10862[5:4] != unexpand_for_this_next_1_case_1_case_0_case_0_case_1;
  assign v0_in_recv_valid = nor_10876 & v0_in_vld;
  assign continuation_9_ctx_4__relative_c_output = sel_10864 == unexpand_for_this_next_1_case_1_case_1_case_0;
  assign __fsm_vvadd_impl_state_17_index = 5'h11;
  assign __for_1_not_exit_state_condition = ~(continuation_9_ctx_4__relative_c_output & ~__for_1_do_break_from_func);
  assign v0_read_pred = 1'h1;
  assign add_10882 = __this_0 + 32'h0000_0001;
  assign __fsm_vvadd_impl_in_state_17 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_17_index;
  assign __fsm_vvadd_impl_go_to_next_state_in_state = ____fsm_vvadd_impl_state_0 == 5'h00 ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h01 ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h02 ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h03 ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h04 ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h05 ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h06 ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h07 ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h08 ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h09 ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h0a ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h0b ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h0c ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h0d ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h0e ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h0f ? v0_read_pred : (____fsm_vvadd_impl_state_0 == 5'h10 ? __for_1_not_exit_state_condition : (____fsm_vvadd_impl_state_0 == 5'h11 ? v0_read_pred : __fsm_vvadd_impl_default_next_state)))))))))))))))));
  assign nand_10891 = ~(~__this_1[0] & ~__this_1[1] & ____fsm_vvadd_impl_state_2);
  assign continuation_4_ctx_3__full_condi_output__2 = (~(continuation_1_ctx_3__full_condi_output__1 & v0_in_recv_valid & eq_10859) ? __this_1 : unexpand_for_this_next_1_case_1_case_1_case_1) == unexpand_for_this_next_1_case_1_case_1_case_1;
  assign continuation_4_ctx_3__full_condi_output = sel_10864 == unexpand_for_this_next_1_case_1_case_1_case_1;
  assign sel_10901 = nand_10891 ? __this_0 : add_10882 & {32{~eq_10859}};
  assign __fsm_vvadd_impl_state_16_index = 5'h10;
  assign and_10936 = continuation_4_ctx_3__full_condi_output__2 & __fsm_vvadd_impl_in_state_0;
  assign nor_10907 = ~(~__fsm_vvadd_impl_in_state_17 | ~__fsm_vvadd_impl_go_to_next_state_in_state | continuation_4_ctx_3__full_condi_output);
  assign eq_10909 = sel_10901 == 32'h0000_000f;
  assign __fsm_vvadd_impl_in_state_16 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_16_index;
  assign v1_in_recv_valid = and_10936 & v1_in_vld;
  assign __fsm_vvadd_impl_state_15_index = 5'h0f;
  assign __fsm_vvadd_impl_state_7_index = 5'h07;
  assign and_10915 = nor_10907 & ~continuation_9_ctx_4__relative_c_output;
  assign and_10917 = __fsm_vvadd_impl_in_state_17 & __fsm_vvadd_impl_go_to_next_state_in_state & continuation_4_ctx_3__full_condi_output;
  assign __for_1_loop_contents_condition = __fsm_vvadd_impl_in_state_16 & continuation_9_ctx_4__relative_c_output;
  assign nor_10933 = ~(continuation_4_ctx_3__full_condi_output | continuation_9_ctx_4__relative_c_output | ~__fsm_vvadd_impl_in_state_17);
  assign and_10968 = continuation_1_ctx_3__full_condi_output__1 & v0_in_recv_valid & __fsm_vvadd_impl_in_state_0;
  assign and_10971 = continuation_4_ctx_3__full_condi_output__2 & v1_in_recv_valid & __fsm_vvadd_impl_in_state_0;
  assign __fsm_vvadd_impl_state_14_index = 5'h0e;
  assign __fsm_vvadd_impl_state_6_index = 5'h06;
  assign __fsm_vvadd_impl_state_13_index = 5'h0d;
  assign __fsm_vvadd_impl_state_5_index = 5'h05;
  assign __fsm_vvadd_impl_in_state_15 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_15_index;
  assign __fsm_vvadd_impl_in_state_7 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_7_index;
  assign __fsm_vvadd_impl_state_11_index = 5'h0b;
  assign __fsm_vvadd_impl_state_3_index = 5'h03;
  assign and_10923 = and_10915 & ~eq_10909;
  assign and_10924 = and_10915 & eq_10909;
  assign and_10925 = and_10917 & ____fsm_vvadd_impl_state_4 & ~eq_10909;
  assign and_10926 = and_10917 & ____fsm_vvadd_impl_state_4 & eq_10909;
  assign and_10927 = and_10917 & ~____fsm_vvadd_impl_state_4 & ~(__this_1[0] | __this_1[1] | ~____fsm_vvadd_impl_state_2);
  assign nor_10928 = ~(~__fsm_vvadd_impl_go_to_next_state_in_state | __fsm_vvadd_impl_in_state_17);
  assign __fsm_vvadd_impl_returns_this_activation_vars = __fsm_vvadd_impl_in_state_17 & __fsm_vvadd_impl_go_to_next_state_in_state;
  assign and_10930 = nor_10907 & continuation_9_ctx_4__relative_c_output;
  assign and_10931 = and_10917 & ~(____fsm_vvadd_impl_state_4 & eq_10909);
  assign p1_all_active_inputs_valid = (~p0___for_1_loop_contents_condition | v0__read_resp_vld) & (~p0___for_1_loop_contents_condition | v1__read_resp_vld) & (~p0_nor_10933 | __c_rd_en__1_delay_reg | __c_ram_zero_latency0_valid_skid_reg) & (~p0_and_10968 | v0__write_completion_vld) & (~p0_and_10971 | v1__write_completion_vld);
  assign p1_all_active_outputs_ready = ~p0_nor_10933 | out_rdy | __out_has_been_sent_reg;
  assign c__read_req_not_pred = ~nor_10933;
  assign c_ram_zero_latency0_from_skid_rdy = ~__c_ram_zero_latency0_valid_skid_reg;
  assign v0__write_req_not_pred = ~and_10968;
  assign v1__write_req_not_pred = ~and_10971;
  assign __fsm_vvadd_impl_state_one = 5'h01;
  assign __fsm_vvadd_impl_state_2_index = 5'h02;
  assign __fsm_vvadd_impl_state_4_index = 5'h04;
  assign __fsm_vvadd_impl_state_8_index = 5'h08;
  assign __fsm_vvadd_impl_state_9_index = 5'h09;
  assign __fsm_vvadd_impl_state_10_index = 5'h0a;
  assign __fsm_vvadd_impl_state_12_index = 5'h0c;
  assign __fsm_vvadd_impl_in_state_14 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_14_index;
  assign __fsm_vvadd_impl_in_state_6 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_6_index;
  assign __fsm_vvadd_impl_in_state_13 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_13_index;
  assign __fsm_vvadd_impl_in_state_5 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_5_index;
  assign and_11053 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_15;
  assign and_11054 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_7;
  assign __fsm_vvadd_impl_in_state_11 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_11_index;
  assign __fsm_vvadd_impl_in_state_3 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_3_index;
  assign __this_0__next_value_predicates = {and_10923, and_10924, and_10925, and_10926, and_10927};
  assign ____fsm_vvadd_impl_state_0__next_value_predicates = {nor_10928, __fsm_vvadd_impl_returns_this_activation_vars};
  assign __this_1__next_value_predicates = {and_10930, and_10926, and_10931, and_10924};
  assign p1_stage_done = p0_valid & p1_all_active_inputs_valid & p1_all_active_outputs_ready;
  assign p1_not_valid = ~p0_valid;
  assign __fsm_vvadd_impl_in_state_1 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_one;
  assign __fsm_vvadd_impl_in_state_2 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_2_index;
  assign __fsm_vvadd_impl_in_state_4 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_4_index;
  assign __fsm_vvadd_impl_in_state_8 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_8_index;
  assign __fsm_vvadd_impl_in_state_9 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_9_index;
  assign __fsm_vvadd_impl_in_state_10 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_10_index;
  assign __fsm_vvadd_impl_in_state_12 = p0_____fsm_vvadd_impl_state_0__1 == __fsm_vvadd_impl_state_12_index;
  assign and_11069 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_14;
  assign and_11070 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_6;
  assign and_11071 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_13;
  assign and_11072 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_5;
  assign or_11074 = and_11053 | and_11054;
  assign and_11075 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_11;
  assign and_11076 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_3;
  assign v0__read_resp_select = p0___for_1_loop_contents_condition ? v0__read_resp : literal_11058;
  assign v1__read_resp_select = p0___for_1_loop_contents_condition ? v1__read_resp : literal_11062;
  assign one_hot_10947 = {__this_0__next_value_predicates[4:0] == 5'h00, __this_0__next_value_predicates[4] && __this_0__next_value_predicates[3:0] == 4'h0, __this_0__next_value_predicates[3] && __this_0__next_value_predicates[2:0] == 3'h0, __this_0__next_value_predicates[2] && __this_0__next_value_predicates[1:0] == 2'h0, __this_0__next_value_predicates[1] && !__this_0__next_value_predicates[0], __this_0__next_value_predicates[0]};
  assign one_hot_10948 = {____fsm_vvadd_impl_state_0__next_value_predicates[1:0] == 2'h0, ____fsm_vvadd_impl_state_0__next_value_predicates[1] && !____fsm_vvadd_impl_state_0__next_value_predicates[0], ____fsm_vvadd_impl_state_0__next_value_predicates[0]};
  assign one_hot_10949 = {__this_1__next_value_predicates[3:0] == 4'h0, __this_1__next_value_predicates[3] && __this_1__next_value_predicates[2:0] == 3'h0, __this_1__next_value_predicates[2] && __this_1__next_value_predicates[1:0] == 2'h0, __this_1__next_value_predicates[1] && !__this_1__next_value_predicates[0], __this_1__next_value_predicates[0]};
  assign p0_enable = p1_stage_done | p1_not_valid;
  assign p0_all_active_outputs_ready = (~__for_1_loop_contents_condition | v0__read_req_rdy | __v0__read_req_has_been_sent_reg) & (~__for_1_loop_contents_condition | v1__read_req_rdy | __v1__read_req_has_been_sent_reg) & (c__read_req_not_pred | c_ram_zero_latency0_from_skid_rdy | __c__read_req_has_been_sent_reg) & (v0__write_req_not_pred | v0__write_req_rdy | __v0__write_req_has_been_sent_reg) & (v1__write_req_not_pred | v1__write_req_rdy | __v1__write_req_has_been_sent_reg);
  assign and_11120 = p0_continuation_9_ctx_4__relative_c_output & p0___fsm_vvadd_impl_in_state_0;
  assign and_11090 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_1;
  assign and_11089 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_2;
  assign and_11087 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_4;
  assign and_11084 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_8;
  assign and_11083 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_9;
  assign and_11082 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_10;
  assign and_11081 = p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_12;
  assign or_11085 = and_11069 | and_11070;
  assign or_11086 = and_11071 | and_11072;
  assign or_11088 = or_11074 | and_11075 | and_11076;
  assign v0_read_response = v0__read_resp_select[31:0];
  assign v1_read_response = v1__read_resp_select[31:0];
  assign c_ram_zero_latency0_select = __c_ram_zero_latency0_valid_skid_reg ? __c_ram_zero_latency0_skid_reg : c_rd_data;
  assign p0_data_enable = p0_enable & p0_all_active_outputs_ready;
  assign __v0__read_req_vld_buf = p0_enable & __for_1_loop_contents_condition;
  assign __v0__read_req_not_has_been_sent = ~__v0__read_req_has_been_sent_reg;
  assign __v1__read_req_not_has_been_sent = ~__v1__read_req_has_been_sent_reg;
  assign __c__read_req_vld_buf = p0_enable & nor_10933;
  assign __c__read_req_not_has_been_sent = ~__c__read_req_has_been_sent_reg;
  assign __v0__write_req_vld_buf = p0_enable & and_10968;
  assign __v0__write_req_not_has_been_sent = ~__v0__write_req_has_been_sent_reg;
  assign __v1__write_req_vld_buf = p0_enable & and_10971;
  assign __v1__write_req_not_has_been_sent = ~__v1__write_req_has_been_sent_reg;
  assign or_11123 = p0___for_1_loop_contents_condition | and_11120 | and_11090 | and_11089 | and_11076 | and_11087 | and_11072 | and_11070 | and_11054 | and_11084 | and_11083 | and_11082 | and_11075 | and_11081 | and_11071 | and_11069 | and_11053;
  assign __out_vld_buf = p1_all_active_inputs_valid & p0_valid & p0_nor_10933;
  assign __out_not_has_been_sent = ~__out_has_been_sent_reg;
  assign and_11437 = p1_stage_done & p0_nor_10933;
  assign v0_write_addr = __this_0[3:0];
  assign c_write_value__16 = v0_read_response + v1_read_response;
  assign and_11395 = and_10923 & p0_data_enable;
  assign and_11396 = and_10924 & p0_data_enable;
  assign and_11397 = and_10925 & p0_data_enable;
  assign and_11398 = and_10926 & p0_data_enable;
  assign and_11399 = and_10927 & p0_data_enable;
  assign and_11406 = nor_10928 & p0_data_enable;
  assign and_11407 = __fsm_vvadd_impl_returns_this_activation_vars & p0_data_enable;
  assign and_11418 = and_10930 & p0_data_enable;
  assign and_11420 = and_10931 & p0_data_enable;
  assign __v0__read_req_valid_and_not_has_been_sent = __v0__read_req_vld_buf & __v0__read_req_not_has_been_sent;
  assign __v1__read_req_valid_and_not_has_been_sent = __v0__read_req_vld_buf & __v1__read_req_not_has_been_sent;
  assign c_rd_en__1 = __c__read_req_vld_buf & __c__read_req_not_has_been_sent;
  assign __v0__write_req_valid_and_not_has_been_sent = __v0__write_req_vld_buf & __v0__write_req_not_has_been_sent;
  assign __v1__write_req_valid_and_not_has_been_sent = __v1__write_req_vld_buf & __v1__write_req_not_has_been_sent;
  assign __c__write_req_vld_buf = p1_all_active_inputs_valid & p0_valid & or_11123;
  assign __c__write_req_not_has_been_sent = ~__c__write_req_has_been_sent_reg;
  assign __out_valid_and_not_has_been_sent = __out_vld_buf & __out_not_has_been_sent;
  assign c_ram_zero_latency0_to_is_not_rdy = ~and_11437;
  assign c_read_addr = nand_10891 ? v0_write_addr : add_10882[3:0];
  assign c__read_resp_select = p0_nor_10933 ? {c_ram_zero_latency0_select} : literal_11126;
  assign v0_read_addr = and_10856[3:0];
  assign v0_in_select = v0_in_recv_valid ? v0_in : 32'h0000_0000;
  assign v1_write_addr = v0_write_addr & {4{~(~__this_1[0] & v0_in_recv_valid)}};
  assign v1_in_select = v1_in_recv_valid ? v1_in : 32'h0000_0000;
  assign __this_0__at_most_one_next_value = and_10923 == one_hot_10947[4] & and_10924 == one_hot_10947[3] & and_10925 == one_hot_10947[2] & and_10926 == one_hot_10947[1] & and_10927 == one_hot_10947[0];
  assign ____fsm_vvadd_impl_state_0__at_most_one_next_value = nor_10928 == one_hot_10948[1] & __fsm_vvadd_impl_returns_this_activation_vars == one_hot_10948[0];
  assign __this_1__at_most_one_next_value = and_10930 == one_hot_10949[3] & and_10926 == one_hot_10949[2] & and_10931 == one_hot_10949[1] & and_10924 == one_hot_10949[0];
  assign concat_11401 = {and_11395, and_11396, and_11397, and_11398, and_11399};
  assign ctx_3__x_literal__1 = 32'h0000_0000;
  assign add_10992 = sel_10901 + 32'h0000_0001;
  assign concat_11409 = {and_11406, and_11407};
  assign __fsm_vvadd_impl_state_plus_one = ____fsm_vvadd_impl_state_0 + __fsm_vvadd_impl_state_one;
  assign concat_11423 = {and_11418, and_11398, and_11420, and_11396};
  assign unexpand_for_this_next_1_case_1_case_0_case_1 = 2'h3;
  assign __for_1_guarded_update_state_elements = ~(~__fsm_vvadd_impl_in_state_16 | ~continuation_9_ctx_4__relative_c_output | and_10856[4]);
  assign __v0__read_req_valid_and_all_active_outputs_ready = __v0__read_req_vld_buf & p0_all_active_outputs_ready;
  assign __v0__read_req_valid_and_ready_txfr = __v0__read_req_valid_and_not_has_been_sent & v0__read_req_rdy;
  assign __v1__read_req_valid_and_ready_txfr = __v1__read_req_valid_and_not_has_been_sent & v1__read_req_rdy;
  assign __c__read_req_valid_and_all_active_outputs_ready = __c__read_req_vld_buf & p0_all_active_outputs_ready;
  assign __c__read_req_valid_and_ready_txfr = c_rd_en__1 & c_ram_zero_latency0_from_skid_rdy;
  assign __v0__write_req_valid_and_all_active_outputs_ready = __v0__write_req_vld_buf & p0_all_active_outputs_ready;
  assign __v0__write_req_valid_and_ready_txfr = __v0__write_req_valid_and_not_has_been_sent & v0__write_req_rdy;
  assign __v1__write_req_valid_and_all_active_outputs_ready = __v1__write_req_vld_buf & p0_all_active_outputs_ready;
  assign __v1__write_req_valid_and_ready_txfr = __v1__write_req_valid_and_not_has_been_sent & v1__write_req_rdy;
  assign __c__write_req_valid_and_all_active_outputs_ready = __c__write_req_vld_buf & p1_all_active_outputs_ready;
  assign c_wr_en__1 = __c__write_req_vld_buf & __c__write_req_not_has_been_sent;
  assign __out_valid_and_all_active_outputs_ready = __out_vld_buf & p1_all_active_outputs_ready;
  assign __out_valid_and_ready_txfr = __out_valid_and_not_has_been_sent & out_rdy;
  assign c_ram_zero_latency0_skid_data_load_en = __c_rd_en__1_delay_reg & c_ram_zero_latency0_from_skid_rdy & c_ram_zero_latency0_to_is_not_rdy;
  assign c_ram_zero_latency0_skid_valid_set_zero = __c_ram_zero_latency0_valid_skid_reg & and_11437;
  assign tuple_10932 = {c_read_addr};
  assign tuple_11122 = {{and_11053 | and_11069 | and_11071 | and_11081 | and_11075 | and_11082 | and_11083 | and_11084 | p0_and_10903, or_11074 | or_11085 | or_11086 | and_11081 | and_11087 | p0_and_10904, or_11088 | or_11085 | and_11082 | and_11089 | p0_and_10905, or_11088 | or_11086 | and_11083 | and_11090 | p0_and_10906}, c_write_value__16 & {32{p0___for_1_loop_contents_condition}}};
  assign c_read_response = c__read_resp_select[31:0];
  assign tuple_10872 = {v0_read_addr};
  assign and_11439 = p1_stage_done & p0___for_1_loop_contents_condition;
  assign or_11572 = ~p0_all_active_outputs_ready | __this_0__at_most_one_next_value | rst;
  assign or_11574 = ~p0_all_active_outputs_ready | ____fsm_vvadd_impl_state_0__at_most_one_next_value | rst;
  assign or_11576 = ~p0_all_active_outputs_ready | __this_1__at_most_one_next_value | rst;
  assign p4_enable = 1'h1;
  assign p3_enable = 1'h1;
  assign p2_enable = 1'h1;
  assign p1_enable = 1'h1;
  assign nand_11132 = ~(p0_continuation_9_ctx_4__relative_c_output & p0___fsm_vvadd_impl_in_state_0);
  assign nand_11133 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_1);
  assign nand_11134 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_2);
  assign nand_11135 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_3);
  assign nand_11136 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_4);
  assign nand_11137 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_5);
  assign nand_11138 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_6);
  assign nand_11139 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_7);
  assign nand_11140 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_8);
  assign nand_11141 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_9);
  assign nand_11142 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_10);
  assign nand_11143 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_11);
  assign nand_11144 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_12);
  assign nand_11145 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_13);
  assign nand_11146 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_14);
  assign nand_11147 = ~(p0_continuation_9_ctx_4__relative_c_output & __fsm_vvadd_impl_in_state_15);
  assign nand_10999 = ~(__fsm_vvadd_impl_in_state_16 & continuation_9_ctx_4__relative_c_output);
  assign and_10903 = __fsm_vvadd_impl_in_state_16 & continuation_9_ctx_4__relative_c_output & and_10856[3];
  assign and_10904 = __fsm_vvadd_impl_in_state_16 & continuation_9_ctx_4__relative_c_output & and_10856[2];
  assign and_10905 = __fsm_vvadd_impl_in_state_16 & continuation_9_ctx_4__relative_c_output & and_10856[1];
  assign and_10906 = __fsm_vvadd_impl_in_state_16 & continuation_9_ctx_4__relative_c_output & and_10856[0];
  assign one_hot_sel_11402 = ctx_3__x_literal__1 & {32{concat_11401[0]}} | ctx_3__x_literal__1 & {32{concat_11401[1]}} | add_10992 & {32{concat_11401[2]}} | ctx_3__x_literal__1 & {32{concat_11401[3]}} | add_10992 & {32{concat_11401[4]}};
  assign or_11403 = and_11395 | and_11396 | and_11397 | and_11398 | and_11399;
  assign one_hot_sel_11410 = __fsm_vvadd_impl_state_0_index & {5{concat_11409[0]}} | __fsm_vvadd_impl_state_plus_one & {5{concat_11409[1]}};
  assign or_11411 = and_11406 | and_11407;
  assign sel_10989 = ____fsm_vvadd_impl_state_0 == 5'h00 ? (____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_valid : ____fsm_vvadd_impl_state_2) : (____fsm_vvadd_impl_state_0 == 5'h01 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h02 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h03 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h04 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h05 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h06 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h07 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h08 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h09 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h0a ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h0b ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h0c ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h0d ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h0e ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h0f ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h10 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 5'h11 ? ____fsm_vvadd_impl_state_2 : __fsm_vvadd_impl_default_next_state)))))))))))))))));
  assign sel_10990 = ____fsm_vvadd_impl_state_0 == 5'h00 ? (____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_valid : ____fsm_vvadd_impl_state_4) : (____fsm_vvadd_impl_state_0 == 5'h01 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h02 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h03 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h04 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h05 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h06 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h07 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h08 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h09 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h0a ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h0b ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h0c ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h0d ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h0e ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h0f ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h10 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 5'h11 ? ____fsm_vvadd_impl_state_4 : __fsm_vvadd_impl_default_next_state)))))))))))))))));
  assign and_11415 = __for_1_loop_contents_condition & p0_data_enable;
  assign one_hot_sel_11424 = unexpand_for_this_next_1_case_1_case_0_case_0_case_1 & {2{concat_11423[0]}} | unexpand_for_this_next_1_case_1_case_1_case_1 & {2{concat_11423[1]}} | unexpand_for_this_next_1_case_1_case_1_case_0 & {2{concat_11423[2]}} | unexpand_for_this_next_1_case_1_case_0_case_1 & {2{concat_11423[3]}};
  assign or_11425 = and_11418 | and_11398 | and_11420 | and_11396;
  assign unexpand_for___for_1_i_next__1_case_1 = add_10862[4:0];
  assign and_11427 = __for_1_guarded_update_state_elements & p0_data_enable;
  assign __v0__read_req_not_stage_load = ~__v0__read_req_valid_and_all_active_outputs_ready;
  assign __v0__read_req_has_been_sent_reg_load_en = __v0__read_req_valid_and_ready_txfr | __v0__read_req_valid_and_all_active_outputs_ready;
  assign __v1__read_req_has_been_sent_reg_load_en = __v1__read_req_valid_and_ready_txfr | __v0__read_req_valid_and_all_active_outputs_ready;
  assign __c__read_req_not_stage_load = ~__c__read_req_valid_and_all_active_outputs_ready;
  assign __c__read_req_has_been_sent_reg_load_en = __c__read_req_valid_and_ready_txfr | __c__read_req_valid_and_all_active_outputs_ready;
  assign __v0__write_req_not_stage_load = ~__v0__write_req_valid_and_all_active_outputs_ready;
  assign __v0__write_req_has_been_sent_reg_load_en = __v0__write_req_valid_and_ready_txfr | __v0__write_req_valid_and_all_active_outputs_ready;
  assign __v1__write_req_not_stage_load = ~__v1__write_req_valid_and_all_active_outputs_ready;
  assign __v1__write_req_has_been_sent_reg_load_en = __v1__write_req_valid_and_ready_txfr | __v1__write_req_valid_and_all_active_outputs_ready;
  assign __c__write_req_not_stage_load = ~__c__write_req_valid_and_all_active_outputs_ready;
  assign __c__write_req_has_been_sent_reg_load_en = c_wr_en__1 | __c__write_req_valid_and_all_active_outputs_ready;
  assign __out_not_stage_load = ~__out_valid_and_all_active_outputs_ready;
  assign __out_has_been_sent_reg_load_en = __out_valid_and_ready_txfr | __out_valid_and_all_active_outputs_ready;
  assign c_ram_zero_latency0_skid_valid_load_en = c_ram_zero_latency0_skid_data_load_en | c_ram_zero_latency0_skid_valid_set_zero;
  always_ff @ (posedge clk) begin
    if (rst) begin
      ____for_1__last_iter_broke <= 1'h1;
      __this_1 <= 2'h0;
      ____for_1_i <= 5'h00;
      __this_0 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_2 <= 1'h0;
      ____fsm_vvadd_impl_state_0 <= 5'h00;
      ____fsm_vvadd_impl_state_4 <= 1'h0;
      ____fsm_vvadd_impl_exited_last_activation <= 1'h1;
      p0_____fsm_vvadd_impl_state_0__1 <= 5'h00;
      p0___fsm_vvadd_impl_in_state_0 <= 1'h0;
      p0_continuation_9_ctx_4__relative_c_output <= 1'h0;
      p0___for_1_loop_contents_condition <= 1'h0;
      p0_nor_10933 <= 1'h0;
      p0_and_10968 <= 1'h0;
      p0_and_10971 <= 1'h0;
      p0_nand_10999 <= 1'h0;
      p0_and_10903 <= 1'h0;
      p0_and_10904 <= 1'h0;
      p0_and_10905 <= 1'h0;
      p0_and_10906 <= 1'h0;
      p1___for_1_loop_contents_condition <= 1'h0;
      p1_and_11120 <= 1'h0;
      p1_and_11090 <= 1'h0;
      p1_and_11089 <= 1'h0;
      p1_and_11076 <= 1'h0;
      p1_and_11087 <= 1'h0;
      p1_and_11072 <= 1'h0;
      p1_and_11070 <= 1'h0;
      p1_and_11054 <= 1'h0;
      p1_and_11084 <= 1'h0;
      p1_and_11083 <= 1'h0;
      p1_and_11082 <= 1'h0;
      p1_and_11075 <= 1'h0;
      p1_and_11081 <= 1'h0;
      p1_and_11071 <= 1'h0;
      p1_and_11069 <= 1'h0;
      p1_and_11053 <= 1'h0;
      p1_or_11123 <= 1'h0;
      p1_nand_10999 <= 1'h0;
      p1_nand_11132 <= 1'h0;
      p1_nand_11133 <= 1'h0;
      p1_nand_11134 <= 1'h0;
      p1_nand_11135 <= 1'h0;
      p1_nand_11136 <= 1'h0;
      p1_nand_11137 <= 1'h0;
      p1_nand_11138 <= 1'h0;
      p1_nand_11139 <= 1'h0;
      p1_nand_11140 <= 1'h0;
      p1_nand_11141 <= 1'h0;
      p1_nand_11142 <= 1'h0;
      p1_nand_11143 <= 1'h0;
      p1_nand_11144 <= 1'h0;
      p1_nand_11145 <= 1'h0;
      p1_nand_11146 <= 1'h0;
      p1_nand_11147 <= 1'h0;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      p4_valid <= 1'h0;
      __v0__read_req_has_been_sent_reg <= 1'h0;
      __v1__read_req_has_been_sent_reg <= 1'h0;
      __c__read_req_has_been_sent_reg <= 1'h0;
      __v0__write_req_has_been_sent_reg <= 1'h0;
      __v1__write_req_has_been_sent_reg <= 1'h0;
      __c__write_req_has_been_sent_reg <= 1'h0;
      __out_has_been_sent_reg <= 1'h0;
      __c_rd_en__1_delay_reg <= 1'h0;
      __c_ram_zero_latency0_skid_reg <= 32'h0000_0000;
      __c_ram_zero_latency0_valid_skid_reg <= 1'h0;
    end else begin
      ____for_1__last_iter_broke <= and_11415 ? __for_1_do_break_from_func : ____for_1__last_iter_broke;
      __this_1 <= or_11425 ? one_hot_sel_11424 : __this_1;
      ____for_1_i <= and_11427 ? unexpand_for___for_1_i_next__1_case_1 : ____for_1_i;
      __this_0 <= or_11403 ? one_hot_sel_11402 : __this_0;
      ____fsm_vvadd_impl_state_2 <= p0_data_enable ? sel_10989 : ____fsm_vvadd_impl_state_2;
      ____fsm_vvadd_impl_state_0 <= or_11411 ? one_hot_sel_11410 : ____fsm_vvadd_impl_state_0;
      ____fsm_vvadd_impl_state_4 <= p0_data_enable ? sel_10990 : ____fsm_vvadd_impl_state_4;
      ____fsm_vvadd_impl_exited_last_activation <= p0_data_enable ? __fsm_vvadd_impl_go_to_next_state_in_state : ____fsm_vvadd_impl_exited_last_activation;
      p0_____fsm_vvadd_impl_state_0__1 <= p0_data_enable ? ____fsm_vvadd_impl_state_0 : p0_____fsm_vvadd_impl_state_0__1;
      p0___fsm_vvadd_impl_in_state_0 <= p0_data_enable ? __fsm_vvadd_impl_in_state_0 : p0___fsm_vvadd_impl_in_state_0;
      p0_continuation_9_ctx_4__relative_c_output <= p0_data_enable ? continuation_9_ctx_4__relative_c_output : p0_continuation_9_ctx_4__relative_c_output;
      p0___for_1_loop_contents_condition <= p0_data_enable ? __for_1_loop_contents_condition : p0___for_1_loop_contents_condition;
      p0_nor_10933 <= p0_data_enable ? nor_10933 : p0_nor_10933;
      p0_and_10968 <= p0_data_enable ? and_10968 : p0_and_10968;
      p0_and_10971 <= p0_data_enable ? and_10971 : p0_and_10971;
      p0_nand_10999 <= p0_data_enable ? nand_10999 : p0_nand_10999;
      p0_and_10903 <= p0_data_enable ? and_10903 : p0_and_10903;
      p0_and_10904 <= p0_data_enable ? and_10904 : p0_and_10904;
      p0_and_10905 <= p0_data_enable ? and_10905 : p0_and_10905;
      p0_and_10906 <= p0_data_enable ? and_10906 : p0_and_10906;
      p1___for_1_loop_contents_condition <= p1_stage_done ? p0___for_1_loop_contents_condition : p1___for_1_loop_contents_condition;
      p1_and_11120 <= p1_stage_done ? and_11120 : p1_and_11120;
      p1_and_11090 <= p1_stage_done ? and_11090 : p1_and_11090;
      p1_and_11089 <= p1_stage_done ? and_11089 : p1_and_11089;
      p1_and_11076 <= p1_stage_done ? and_11076 : p1_and_11076;
      p1_and_11087 <= p1_stage_done ? and_11087 : p1_and_11087;
      p1_and_11072 <= p1_stage_done ? and_11072 : p1_and_11072;
      p1_and_11070 <= p1_stage_done ? and_11070 : p1_and_11070;
      p1_and_11054 <= p1_stage_done ? and_11054 : p1_and_11054;
      p1_and_11084 <= p1_stage_done ? and_11084 : p1_and_11084;
      p1_and_11083 <= p1_stage_done ? and_11083 : p1_and_11083;
      p1_and_11082 <= p1_stage_done ? and_11082 : p1_and_11082;
      p1_and_11075 <= p1_stage_done ? and_11075 : p1_and_11075;
      p1_and_11081 <= p1_stage_done ? and_11081 : p1_and_11081;
      p1_and_11071 <= p1_stage_done ? and_11071 : p1_and_11071;
      p1_and_11069 <= p1_stage_done ? and_11069 : p1_and_11069;
      p1_and_11053 <= p1_stage_done ? and_11053 : p1_and_11053;
      p1_or_11123 <= p1_stage_done ? or_11123 : p1_or_11123;
      p1_nand_10999 <= p1_stage_done ? p0_nand_10999 : p1_nand_10999;
      p1_nand_11132 <= p1_stage_done ? nand_11132 : p1_nand_11132;
      p1_nand_11133 <= p1_stage_done ? nand_11133 : p1_nand_11133;
      p1_nand_11134 <= p1_stage_done ? nand_11134 : p1_nand_11134;
      p1_nand_11135 <= p1_stage_done ? nand_11135 : p1_nand_11135;
      p1_nand_11136 <= p1_stage_done ? nand_11136 : p1_nand_11136;
      p1_nand_11137 <= p1_stage_done ? nand_11137 : p1_nand_11137;
      p1_nand_11138 <= p1_stage_done ? nand_11138 : p1_nand_11138;
      p1_nand_11139 <= p1_stage_done ? nand_11139 : p1_nand_11139;
      p1_nand_11140 <= p1_stage_done ? nand_11140 : p1_nand_11140;
      p1_nand_11141 <= p1_stage_done ? nand_11141 : p1_nand_11141;
      p1_nand_11142 <= p1_stage_done ? nand_11142 : p1_nand_11142;
      p1_nand_11143 <= p1_stage_done ? nand_11143 : p1_nand_11143;
      p1_nand_11144 <= p1_stage_done ? nand_11144 : p1_nand_11144;
      p1_nand_11145 <= p1_stage_done ? nand_11145 : p1_nand_11145;
      p1_nand_11146 <= p1_stage_done ? nand_11146 : p1_nand_11146;
      p1_nand_11147 <= p1_stage_done ? nand_11147 : p1_nand_11147;
      p0_valid <= p0_enable ? p0_all_active_outputs_ready : p0_valid;
      p1_valid <= p1_enable ? p1_stage_done : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      p4_valid <= p4_enable ? p3_valid : p4_valid;
      __v0__read_req_has_been_sent_reg <= __v0__read_req_has_been_sent_reg_load_en ? __v0__read_req_not_stage_load : __v0__read_req_has_been_sent_reg;
      __v1__read_req_has_been_sent_reg <= __v1__read_req_has_been_sent_reg_load_en ? __v0__read_req_not_stage_load : __v1__read_req_has_been_sent_reg;
      __c__read_req_has_been_sent_reg <= __c__read_req_has_been_sent_reg_load_en ? __c__read_req_not_stage_load : __c__read_req_has_been_sent_reg;
      __v0__write_req_has_been_sent_reg <= __v0__write_req_has_been_sent_reg_load_en ? __v0__write_req_not_stage_load : __v0__write_req_has_been_sent_reg;
      __v1__write_req_has_been_sent_reg <= __v1__write_req_has_been_sent_reg_load_en ? __v1__write_req_not_stage_load : __v1__write_req_has_been_sent_reg;
      __c__write_req_has_been_sent_reg <= __c__write_req_has_been_sent_reg_load_en ? __c__write_req_not_stage_load : __c__write_req_has_been_sent_reg;
      __out_has_been_sent_reg <= __out_has_been_sent_reg_load_en ? __out_not_stage_load : __out_has_been_sent_reg;
      __c_rd_en__1_delay_reg <= c_rd_en__1;
      __c_ram_zero_latency0_skid_reg <= c_ram_zero_latency0_skid_data_load_en ? c_rd_data : __c_ram_zero_latency0_skid_reg;
      __c_ram_zero_latency0_valid_skid_reg <= c_ram_zero_latency0_skid_valid_load_en ? c_ram_zero_latency0_from_skid_rdy : __c_ram_zero_latency0_valid_skid_reg;
    end
  end
  assign out = c_read_response;
  assign out_vld = __out_valid_and_not_has_been_sent;
  assign v0__read_req = tuple_10872;
  assign v0__read_req_vld = __v0__read_req_valid_and_not_has_been_sent;
  assign v0__read_resp_rdy = and_11439;
  assign v0__write_completion_rdy = p1_stage_done & p0_and_10968;
  assign v0__write_req = {v0_write_addr, v0_in_select};
  assign v0__write_req_vld = __v0__write_req_valid_and_not_has_been_sent;
  assign v0_in_rdy = p0_data_enable & nor_10876;
  assign v1__read_req = tuple_10872;
  assign v1__read_req_vld = __v1__read_req_valid_and_not_has_been_sent;
  assign v1__read_resp_rdy = and_11439;
  assign v1__write_completion_rdy = p1_stage_done & p0_and_10971;
  assign v1__write_req = {v1_write_addr, v1_in_select};
  assign v1__write_req_vld = __v1__write_req_valid_and_not_has_been_sent;
  assign v1_in_rdy = p0_data_enable & and_10936;
  assign c_rd_addr = tuple_10932[3:0];
  assign c_rd_en = c_rd_en__1;
  assign c_wr_addr = tuple_11122[35:32];
  assign c_wr_data = tuple_11122[31:0];
  assign c_wr_en = c_wr_en__1;
  `ifdef ASSERT_ON
  __this_0__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_11572))) or_11572) else $fatal(0, "More than one next_value fired for state element: this_0");
  ____fsm_vvadd_impl_state_0__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_11574))) or_11574) else $fatal(0, "More than one next_value fired for state element: __fsm_vvadd_impl_state_0");
  __this_1__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_11576))) or_11576) else $fatal(0, "More than one next_value fired for state element: this_1");
  `endif  // ASSERT_ON
endmodule
