module xls_vvadd(
  input wire clk,
  input wire rst,
  input wire out_rdy,
  input wire [31:0] v0_in,
  input wire v0_in_vld,
  input wire [31:0] v1_in,
  input wire v1_in_vld,
  output wire [31:0] out,
  output wire out_vld,
  output wire v0_in_rdy,
  output wire v1_in_rdy
);
  wire [31:0] ____for_1_c_init[16];
  assign ____for_1_c_init = '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000};
  wire [31:0] literal_22756[16];
  assign literal_22756 = '{32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000, 32'h0000_0000};
  reg ____for_1__last_iter_broke;
  reg [5:0] ____fsm_vvadd_impl_state_0;
  reg [4:0] ____for_1_i;
  reg ____fsm_vvadd_impl_exited_last_activation;
  reg [31:0] ____fsm_vvadd_impl_state_32;
  reg [31:0] ____fsm_vvadd_impl_state_1;
  reg [31:0] ____fsm_vvadd_impl_state_2;
  reg [31:0] ____fsm_vvadd_impl_state_3;
  reg [31:0] ____fsm_vvadd_impl_state_4;
  reg [31:0] ____fsm_vvadd_impl_state_5;
  reg [31:0] ____fsm_vvadd_impl_state_6;
  reg [31:0] ____fsm_vvadd_impl_state_7;
  reg [31:0] ____fsm_vvadd_impl_state_8;
  reg [31:0] ____fsm_vvadd_impl_state_9;
  reg [31:0] ____fsm_vvadd_impl_state_10;
  reg [31:0] ____fsm_vvadd_impl_state_11;
  reg [31:0] ____fsm_vvadd_impl_state_12;
  reg [31:0] ____fsm_vvadd_impl_state_13;
  reg [31:0] ____fsm_vvadd_impl_state_14;
  reg [31:0] ____fsm_vvadd_impl_state_15;
  reg [31:0] ____fsm_vvadd_impl_state_16;
  reg [31:0] ____fsm_vvadd_impl_state_17;
  reg [31:0] ____fsm_vvadd_impl_state_18;
  reg [31:0] ____fsm_vvadd_impl_state_19;
  reg [31:0] ____fsm_vvadd_impl_state_20;
  reg [31:0] ____fsm_vvadd_impl_state_21;
  reg [31:0] ____fsm_vvadd_impl_state_22;
  reg [31:0] ____fsm_vvadd_impl_state_23;
  reg [31:0] ____fsm_vvadd_impl_state_24;
  reg [31:0] ____fsm_vvadd_impl_state_25;
  reg [31:0] ____fsm_vvadd_impl_state_26;
  reg [31:0] ____fsm_vvadd_impl_state_27;
  reg [31:0] ____fsm_vvadd_impl_state_28;
  reg [31:0] ____fsm_vvadd_impl_state_29;
  reg [31:0] ____fsm_vvadd_impl_state_30;
  reg [31:0] ____fsm_vvadd_impl_state_31;
  reg [31:0] ____for_1_c[16];
  wire __fsm_vvadd_impl_default_next_state;
  wire [4:0] and_22811;
  wire [5:0] __fsm_vvadd_impl_state_1_index;
  wire [5:0] __fsm_vvadd_impl_state_30_index;
  wire [5:0] add_22847;
  wire [5:0] __fsm_vvadd_impl_state_15_index;
  wire [5:0] __fsm_vvadd_impl_state_16_index;
  wire [5:0] __fsm_vvadd_impl_state_17_index;
  wire [5:0] __fsm_vvadd_impl_state_18_index;
  wire [5:0] __fsm_vvadd_impl_state_19_index;
  wire [5:0] __fsm_vvadd_impl_state_20_index;
  wire [5:0] __fsm_vvadd_impl_state_21_index;
  wire [5:0] __fsm_vvadd_impl_state_22_index;
  wire [5:0] __fsm_vvadd_impl_state_23_index;
  wire [5:0] __fsm_vvadd_impl_state_24_index;
  wire [5:0] __fsm_vvadd_impl_state_25_index;
  wire [5:0] __fsm_vvadd_impl_state_26_index;
  wire [5:0] __fsm_vvadd_impl_state_27_index;
  wire [5:0] __fsm_vvadd_impl_state_28_index;
  wire [5:0] __fsm_vvadd_impl_state_29_index;
  wire __fsm_vvadd_impl_in_state_30;
  wire __fsm_vvadd_impl_in_state_15;
  wire __fsm_vvadd_impl_in_state_16;
  wire __fsm_vvadd_impl_in_state_17;
  wire __fsm_vvadd_impl_in_state_18;
  wire __fsm_vvadd_impl_in_state_19;
  wire __fsm_vvadd_impl_in_state_20;
  wire __fsm_vvadd_impl_in_state_21;
  wire __fsm_vvadd_impl_in_state_22;
  wire __fsm_vvadd_impl_in_state_23;
  wire __fsm_vvadd_impl_in_state_24;
  wire __fsm_vvadd_impl_in_state_25;
  wire __fsm_vvadd_impl_in_state_26;
  wire __fsm_vvadd_impl_in_state_27;
  wire __fsm_vvadd_impl_in_state_28;
  wire __fsm_vvadd_impl_in_state_29;
  wire and_22843;
  wire __for_1_do_break_from_func;
  wire continuation_1_literal;
  wire or_22846;
  wire __fsm_vvadd_impl_go_to_next_state_in_state;
  wire [5:0] __fsm_vvadd_impl_final_state_index;
  wire [5:0] __fsm_vvadd_impl_state_31_index;
  wire [5:0] __fsm_vvadd_impl_state_32_index;
  wire [5:0] __fsm_vvadd_impl_state_33_index;
  wire [5:0] __fsm_vvadd_impl_state_34_index;
  wire [5:0] __fsm_vvadd_impl_state_35_index;
  wire [5:0] __fsm_vvadd_impl_state_36_index;
  wire [5:0] __fsm_vvadd_impl_state_37_index;
  wire [5:0] __fsm_vvadd_impl_state_38_index;
  wire [5:0] __fsm_vvadd_impl_state_39_index;
  wire [5:0] __fsm_vvadd_impl_state_40_index;
  wire [5:0] __fsm_vvadd_impl_state_41_index;
  wire [5:0] __fsm_vvadd_impl_state_42_index;
  wire [5:0] __fsm_vvadd_impl_state_43_index;
  wire [5:0] __fsm_vvadd_impl_state_44_index;
  wire [31:0] v1_in_select;
  wire __fsm_vvadd_impl_in_final_state;
  wire nor_22913;
  wire and_22972;
  wire __fsm_vvadd_impl_in_state_31;
  wire __fsm_vvadd_impl_in_state_32;
  wire __fsm_vvadd_impl_in_state_33;
  wire __fsm_vvadd_impl_in_state_34;
  wire __fsm_vvadd_impl_in_state_35;
  wire __fsm_vvadd_impl_in_state_36;
  wire __fsm_vvadd_impl_in_state_37;
  wire __fsm_vvadd_impl_in_state_38;
  wire __fsm_vvadd_impl_in_state_39;
  wire __fsm_vvadd_impl_in_state_40;
  wire __fsm_vvadd_impl_in_state_41;
  wire __fsm_vvadd_impl_in_state_42;
  wire __fsm_vvadd_impl_in_state_43;
  wire __fsm_vvadd_impl_in_state_44;
  wire [26:0] leading_bits___for_1_i;
  wire [31:0] v1_in_recv_value__15;
  wire nor_22917;
  wire and_22918;
  wire v1_in_not_pred;
  wire v0_in_not_pred;
  wire or_23090;
  wire [31:0] concat_22877;
  wire [31:0] __fsm_vvadd_impl_state_30_select_v1_in_recv_before_loop;
  wire [1:0] ____fsm_vvadd_impl_state_0__next_value_predicates;
  wire out_not_pred;
  wire [5:0] __fsm_vvadd_impl_state_0_index;
  wire [5:0] __fsm_vvadd_impl_state_2_index;
  wire [5:0] __fsm_vvadd_impl_state_3_index;
  wire [5:0] __fsm_vvadd_impl_state_4_index;
  wire [5:0] __fsm_vvadd_impl_state_5_index;
  wire [5:0] __fsm_vvadd_impl_state_6_index;
  wire [5:0] __fsm_vvadd_impl_state_7_index;
  wire [5:0] __fsm_vvadd_impl_state_8_index;
  wire [5:0] __fsm_vvadd_impl_state_9_index;
  wire [5:0] __fsm_vvadd_impl_state_10_index;
  wire [5:0] __fsm_vvadd_impl_state_11_index;
  wire [5:0] __fsm_vvadd_impl_state_12_index;
  wire [5:0] __fsm_vvadd_impl_state_13_index;
  wire [5:0] __fsm_vvadd_impl_state_14_index;
  wire [2:0] one_hot_22988;
  wire p0_all_active_inputs_valid;
  wire __fsm_vvadd_impl_in_state_0;
  wire __fsm_vvadd_impl_in_state_1;
  wire __fsm_vvadd_impl_in_state_2;
  wire __fsm_vvadd_impl_in_state_3;
  wire __fsm_vvadd_impl_in_state_4;
  wire __fsm_vvadd_impl_in_state_5;
  wire __fsm_vvadd_impl_in_state_6;
  wire __fsm_vvadd_impl_in_state_7;
  wire __fsm_vvadd_impl_in_state_8;
  wire __fsm_vvadd_impl_in_state_9;
  wire __fsm_vvadd_impl_in_state_10;
  wire __fsm_vvadd_impl_in_state_11;
  wire __fsm_vvadd_impl_in_state_12;
  wire __fsm_vvadd_impl_in_state_13;
  wire __fsm_vvadd_impl_in_state_14;
  wire [31:0] sel_22938[16];
  wire [31:0] add_22939;
  wire p0_stage_done;
  wire [31:0] v0_in_select;
  wire [31:0] sign_ext_22957;
  wire [31:0] array_update_22987[16];
  wire [31:0] v0_in_recv_value;
  wire [31:0] v0_in_recv_value__1;
  wire [31:0] v0_in_recv_value__2;
  wire [31:0] v0_in_recv_value__3;
  wire [31:0] v0_in_recv_value__4;
  wire [31:0] v0_in_recv_value__5;
  wire [31:0] v0_in_recv_value__6;
  wire [31:0] v0_in_recv_value__7;
  wire [31:0] v0_in_recv_value__8;
  wire [31:0] v0_in_recv_value__9;
  wire [31:0] v0_in_recv_value__10;
  wire [31:0] v0_in_recv_value__11;
  wire [31:0] v0_in_recv_value__12;
  wire [31:0] v0_in_recv_value__13;
  wire [31:0] v0_in_recv_value__14;
  wire [31:0] v0_in_recv_value__15;
  wire [31:0] v1_in_recv_value;
  wire [31:0] v1_in_recv_value__1;
  wire [31:0] v1_in_recv_value__2;
  wire [31:0] v1_in_recv_value__3;
  wire [31:0] v1_in_recv_value__4;
  wire [31:0] v1_in_recv_value__5;
  wire [31:0] v1_in_recv_value__6;
  wire [31:0] v1_in_recv_value__7;
  wire [31:0] v1_in_recv_value__8;
  wire [31:0] v1_in_recv_value__9;
  wire [31:0] v1_in_recv_value__10;
  wire [31:0] v1_in_recv_value__11;
  wire [31:0] v1_in_recv_value__12;
  wire [31:0] v1_in_recv_value__13;
  wire [31:0] v1_in_recv_value__14;
  wire [15:0] concat_23037;
  wire [31:0] out_send_value__15;
  wire [31:0] out_send_value__14;
  wire [31:0] out_send_value__13;
  wire [31:0] out_send_value__12;
  wire [31:0] out_send_value__11;
  wire [31:0] out_send_value__10;
  wire [31:0] out_send_value__9;
  wire [31:0] out_send_value__8;
  wire [31:0] out_send_value__7;
  wire [31:0] out_send_value__6;
  wire [31:0] out_send_value__5;
  wire [31:0] out_send_value__4;
  wire [31:0] out_send_value__3;
  wire [31:0] out_send_value__2;
  wire [31:0] out_send_value__1;
  wire [31:0] out_send_value;
  wire ____fsm_vvadd_impl_state_0__at_most_one_next_value;
  wire [1:0] concat_23234;
  wire [5:0] __fsm_vvadd_impl_state_plus_one;
  wire [31:0] __fsm_vvadd_impl_state_0_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_1_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_2_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_3_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_4_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_5_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_6_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_7_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_8_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_9_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_10_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_11_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_12_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_13_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_14_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_15_select_v0_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_15_select_v1_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_16_select_v1_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_17_select_v1_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_18_select_v1_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_19_select_v1_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_20_select_v1_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_21_select_v1_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_22_select_v1_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_23_select_v1_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_24_select_v1_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_25_select_v1_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_26_select_v1_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_27_select_v1_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_28_select_v1_in_recv_before_loop;
  wire [31:0] __fsm_vvadd_impl_state_29_select_v1_in_recv_before_loop;
  wire __for_1_guarded_update_state_elements;
  wire or_23326;
  wire [5:0] one_hot_sel_23235;
  wire and_23283;
  wire [31:0] sel_23095;
  wire [31:0] sel_23096;
  wire [31:0] sel_23097;
  wire [31:0] sel_23098;
  wire [31:0] sel_23099;
  wire [31:0] sel_23100;
  wire [31:0] sel_23101;
  wire [31:0] sel_23102;
  wire [31:0] sel_23103;
  wire [31:0] sel_23104;
  wire [31:0] sel_23105;
  wire [31:0] sel_23106;
  wire [31:0] sel_23107;
  wire [31:0] sel_23108;
  wire [31:0] sel_23109;
  wire [31:0] sel_23110;
  wire [31:0] sel_23111;
  wire [31:0] sel_23112;
  wire [31:0] sel_23113;
  wire [31:0] sel_23114;
  wire [31:0] sel_23115;
  wire [31:0] sel_23116;
  wire [31:0] sel_23117;
  wire [31:0] sel_23118;
  wire [31:0] sel_23119;
  wire [31:0] sel_23120;
  wire [31:0] sel_23121;
  wire [31:0] sel_23122;
  wire [31:0] sel_23123;
  wire [31:0] sel_23124;
  wire [31:0] sel_23125;
  wire [31:0] sel_23126;
  wire and_23317;
  wire and_23319;
  wire [4:0] unexpand_for___for_1_i_next__1_case_1;
  assign __fsm_vvadd_impl_default_next_state = 1'h0;
  assign and_22811 = {5{~____for_1__last_iter_broke}} & ____for_1_i;
  assign __fsm_vvadd_impl_state_1_index = 6'h01;
  assign __fsm_vvadd_impl_state_30_index = 6'h1e;
  assign add_22847 = {__fsm_vvadd_impl_default_next_state, and_22811} + __fsm_vvadd_impl_state_1_index;
  assign __fsm_vvadd_impl_state_15_index = 6'h0f;
  assign __fsm_vvadd_impl_state_16_index = 6'h10;
  assign __fsm_vvadd_impl_state_17_index = 6'h11;
  assign __fsm_vvadd_impl_state_18_index = 6'h12;
  assign __fsm_vvadd_impl_state_19_index = 6'h13;
  assign __fsm_vvadd_impl_state_20_index = 6'h14;
  assign __fsm_vvadd_impl_state_21_index = 6'h15;
  assign __fsm_vvadd_impl_state_22_index = 6'h16;
  assign __fsm_vvadd_impl_state_23_index = 6'h17;
  assign __fsm_vvadd_impl_state_24_index = 6'h18;
  assign __fsm_vvadd_impl_state_25_index = 6'h19;
  assign __fsm_vvadd_impl_state_26_index = 6'h1a;
  assign __fsm_vvadd_impl_state_27_index = 6'h1b;
  assign __fsm_vvadd_impl_state_28_index = 6'h1c;
  assign __fsm_vvadd_impl_state_29_index = 6'h1d;
  assign __fsm_vvadd_impl_in_state_30 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_30_index;
  assign __fsm_vvadd_impl_in_state_15 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_15_index;
  assign __fsm_vvadd_impl_in_state_16 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_16_index;
  assign __fsm_vvadd_impl_in_state_17 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_17_index;
  assign __fsm_vvadd_impl_in_state_18 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_18_index;
  assign __fsm_vvadd_impl_in_state_19 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_19_index;
  assign __fsm_vvadd_impl_in_state_20 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_20_index;
  assign __fsm_vvadd_impl_in_state_21 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_21_index;
  assign __fsm_vvadd_impl_in_state_22 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_22_index;
  assign __fsm_vvadd_impl_in_state_23 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_23_index;
  assign __fsm_vvadd_impl_in_state_24 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_24_index;
  assign __fsm_vvadd_impl_in_state_25 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_25_index;
  assign __fsm_vvadd_impl_in_state_26 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_26_index;
  assign __fsm_vvadd_impl_in_state_27 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_27_index;
  assign __fsm_vvadd_impl_in_state_28 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_28_index;
  assign __fsm_vvadd_impl_in_state_29 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_29_index;
  assign and_22843 = ____for_1__last_iter_broke & ____fsm_vvadd_impl_exited_last_activation & __fsm_vvadd_impl_in_state_30;
  assign __for_1_do_break_from_func = add_22847[5:4] != 2'h0;
  assign continuation_1_literal = 1'h1;
  assign or_22846 = __fsm_vvadd_impl_in_state_15 | __fsm_vvadd_impl_in_state_16 | __fsm_vvadd_impl_in_state_17 | __fsm_vvadd_impl_in_state_18 | __fsm_vvadd_impl_in_state_19 | __fsm_vvadd_impl_in_state_20 | __fsm_vvadd_impl_in_state_21 | __fsm_vvadd_impl_in_state_22 | __fsm_vvadd_impl_in_state_23 | __fsm_vvadd_impl_in_state_24 | __fsm_vvadd_impl_in_state_25 | __fsm_vvadd_impl_in_state_26 | __fsm_vvadd_impl_in_state_27 | __fsm_vvadd_impl_in_state_28 | __fsm_vvadd_impl_in_state_29 | and_22843;
  assign __fsm_vvadd_impl_go_to_next_state_in_state = ____fsm_vvadd_impl_state_0 == 6'h00 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h01 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h02 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h03 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h04 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h05 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h06 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h07 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h08 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h09 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h0a ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h0b ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h0c ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h0d ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h0e ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h0f ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h10 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h11 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h12 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h13 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h14 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h15 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h16 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h17 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h18 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h19 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h1a ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h1b ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h1c ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h1d ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h1e ? __for_1_do_break_from_func : (____fsm_vvadd_impl_state_0 == 6'h1f ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h20 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h21 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h22 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h23 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h24 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h25 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h26 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h27 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h28 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h29 ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h2a ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h2b ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h2c ? continuation_1_literal : (____fsm_vvadd_impl_state_0 == 6'h2d ? continuation_1_literal : __fsm_vvadd_impl_default_next_state)))))))))))))))))))))))))))))))))))))))))))));
  assign __fsm_vvadd_impl_final_state_index = 6'h2d;
  assign __fsm_vvadd_impl_state_31_index = 6'h1f;
  assign __fsm_vvadd_impl_state_32_index = 6'h20;
  assign __fsm_vvadd_impl_state_33_index = 6'h21;
  assign __fsm_vvadd_impl_state_34_index = 6'h22;
  assign __fsm_vvadd_impl_state_35_index = 6'h23;
  assign __fsm_vvadd_impl_state_36_index = 6'h24;
  assign __fsm_vvadd_impl_state_37_index = 6'h25;
  assign __fsm_vvadd_impl_state_38_index = 6'h26;
  assign __fsm_vvadd_impl_state_39_index = 6'h27;
  assign __fsm_vvadd_impl_state_40_index = 6'h28;
  assign __fsm_vvadd_impl_state_41_index = 6'h29;
  assign __fsm_vvadd_impl_state_42_index = 6'h2a;
  assign __fsm_vvadd_impl_state_43_index = 6'h2b;
  assign __fsm_vvadd_impl_state_44_index = 6'h2c;
  assign v1_in_select = or_22846 ? v1_in : 32'h0000_0000;
  assign __fsm_vvadd_impl_in_final_state = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_final_state_index;
  assign nor_22913 = ~(____fsm_vvadd_impl_state_0[4] | ____fsm_vvadd_impl_state_0[5]);
  assign and_22972 = __for_1_do_break_from_func & __fsm_vvadd_impl_in_state_30;
  assign __fsm_vvadd_impl_in_state_31 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_31_index;
  assign __fsm_vvadd_impl_in_state_32 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_32_index;
  assign __fsm_vvadd_impl_in_state_33 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_33_index;
  assign __fsm_vvadd_impl_in_state_34 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_34_index;
  assign __fsm_vvadd_impl_in_state_35 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_35_index;
  assign __fsm_vvadd_impl_in_state_36 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_36_index;
  assign __fsm_vvadd_impl_in_state_37 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_37_index;
  assign __fsm_vvadd_impl_in_state_38 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_38_index;
  assign __fsm_vvadd_impl_in_state_39 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_39_index;
  assign __fsm_vvadd_impl_in_state_40 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_40_index;
  assign __fsm_vvadd_impl_in_state_41 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_41_index;
  assign __fsm_vvadd_impl_in_state_42 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_42_index;
  assign __fsm_vvadd_impl_in_state_43 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_43_index;
  assign __fsm_vvadd_impl_in_state_44 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_44_index;
  assign leading_bits___for_1_i = 27'h000_0000;
  assign v1_in_recv_value__15 = v1_in_select & {32{and_22843}};
  assign nor_22917 = ~(~__fsm_vvadd_impl_go_to_next_state_in_state | __fsm_vvadd_impl_in_final_state);
  assign and_22918 = __fsm_vvadd_impl_go_to_next_state_in_state & __fsm_vvadd_impl_in_final_state;
  assign v1_in_not_pred = ~or_22846;
  assign v0_in_not_pred = ~nor_22913;
  assign or_23090 = and_22972 | __fsm_vvadd_impl_in_state_31 | __fsm_vvadd_impl_in_state_32 | __fsm_vvadd_impl_in_state_33 | __fsm_vvadd_impl_in_state_34 | __fsm_vvadd_impl_in_state_35 | __fsm_vvadd_impl_in_state_36 | __fsm_vvadd_impl_in_state_37 | __fsm_vvadd_impl_in_state_38 | __fsm_vvadd_impl_in_state_39 | __fsm_vvadd_impl_in_state_40 | __fsm_vvadd_impl_in_state_41 | __fsm_vvadd_impl_in_state_42 | __fsm_vvadd_impl_in_state_43 | __fsm_vvadd_impl_in_state_44 | __fsm_vvadd_impl_in_final_state;
  assign concat_22877 = {leading_bits___for_1_i, and_22811};
  assign __fsm_vvadd_impl_state_30_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__15 : ____fsm_vvadd_impl_state_32;
  assign ____fsm_vvadd_impl_state_0__next_value_predicates = {nor_22917, and_22918};
  assign out_not_pred = ~or_23090;
  assign __fsm_vvadd_impl_state_0_index = 6'h00;
  assign __fsm_vvadd_impl_state_2_index = 6'h02;
  assign __fsm_vvadd_impl_state_3_index = 6'h03;
  assign __fsm_vvadd_impl_state_4_index = 6'h04;
  assign __fsm_vvadd_impl_state_5_index = 6'h05;
  assign __fsm_vvadd_impl_state_6_index = 6'h06;
  assign __fsm_vvadd_impl_state_7_index = 6'h07;
  assign __fsm_vvadd_impl_state_8_index = 6'h08;
  assign __fsm_vvadd_impl_state_9_index = 6'h09;
  assign __fsm_vvadd_impl_state_10_index = 6'h0a;
  assign __fsm_vvadd_impl_state_11_index = 6'h0b;
  assign __fsm_vvadd_impl_state_12_index = 6'h0c;
  assign __fsm_vvadd_impl_state_13_index = 6'h0d;
  assign __fsm_vvadd_impl_state_14_index = 6'h0e;
  assign one_hot_22988 = {____fsm_vvadd_impl_state_0__next_value_predicates[1:0] == 2'h0, ____fsm_vvadd_impl_state_0__next_value_predicates[1] && !____fsm_vvadd_impl_state_0__next_value_predicates[0], ____fsm_vvadd_impl_state_0__next_value_predicates[0]};
  assign p0_all_active_inputs_valid = (v1_in_not_pred | v1_in_vld) & (v0_in_not_pred | v0_in_vld);
  assign __fsm_vvadd_impl_in_state_0 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_0_index;
  assign __fsm_vvadd_impl_in_state_1 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_1_index;
  assign __fsm_vvadd_impl_in_state_2 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_2_index;
  assign __fsm_vvadd_impl_in_state_3 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_3_index;
  assign __fsm_vvadd_impl_in_state_4 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_4_index;
  assign __fsm_vvadd_impl_in_state_5 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_5_index;
  assign __fsm_vvadd_impl_in_state_6 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_6_index;
  assign __fsm_vvadd_impl_in_state_7 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_7_index;
  assign __fsm_vvadd_impl_in_state_8 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_8_index;
  assign __fsm_vvadd_impl_in_state_9 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_9_index;
  assign __fsm_vvadd_impl_in_state_10 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_10_index;
  assign __fsm_vvadd_impl_in_state_11 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_11_index;
  assign __fsm_vvadd_impl_in_state_12 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_12_index;
  assign __fsm_vvadd_impl_in_state_13 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_13_index;
  assign __fsm_vvadd_impl_in_state_14 = ____fsm_vvadd_impl_state_0 == __fsm_vvadd_impl_state_14_index;
  assign sel_22938 = ____for_1__last_iter_broke == 1'h0 ? ____for_1_c : literal_22756;
  assign add_22939 = (concat_22877 == 32'h0000_0000 ? ____fsm_vvadd_impl_state_1 : (concat_22877 == 32'h0000_0001 ? ____fsm_vvadd_impl_state_2 : (concat_22877 == 32'h0000_0002 ? ____fsm_vvadd_impl_state_3 : (concat_22877 == 32'h0000_0003 ? ____fsm_vvadd_impl_state_4 : (concat_22877 == 32'h0000_0004 ? ____fsm_vvadd_impl_state_5 : (concat_22877 == 32'h0000_0005 ? ____fsm_vvadd_impl_state_6 : (concat_22877 == 32'h0000_0006 ? ____fsm_vvadd_impl_state_7 : (concat_22877 == 32'h0000_0007 ? ____fsm_vvadd_impl_state_8 : (concat_22877 == 32'h0000_0008 ? ____fsm_vvadd_impl_state_9 : (concat_22877 == 32'h0000_0009 ? ____fsm_vvadd_impl_state_10 : (concat_22877 == 32'h0000_000a ? ____fsm_vvadd_impl_state_11 : (concat_22877 == 32'h0000_000b ? ____fsm_vvadd_impl_state_12 : (concat_22877 == 32'h0000_000c ? ____fsm_vvadd_impl_state_13 : (concat_22877 == 32'h0000_000d ? ____fsm_vvadd_impl_state_14 : (concat_22877 == 32'h0000_000e ? ____fsm_vvadd_impl_state_15 : ____fsm_vvadd_impl_state_16))))))))))))))) + (concat_22877 == 32'h0000_0000 ? ____fsm_vvadd_impl_state_17 : (concat_22877 == 32'h0000_0001 ? ____fsm_vvadd_impl_state_18 : (concat_22877 == 32'h0000_0002 ? ____fsm_vvadd_impl_state_19 : (concat_22877 == 32'h0000_0003 ? ____fsm_vvadd_impl_state_20 : (concat_22877 == 32'h0000_0004 ? ____fsm_vvadd_impl_state_21 : (concat_22877 == 32'h0000_0005 ? ____fsm_vvadd_impl_state_22 : (concat_22877 == 32'h0000_0006 ? ____fsm_vvadd_impl_state_23 : (concat_22877 == 32'h0000_0007 ? ____fsm_vvadd_impl_state_24 : (concat_22877 == 32'h0000_0008 ? ____fsm_vvadd_impl_state_25 : (concat_22877 == 32'h0000_0009 ? ____fsm_vvadd_impl_state_26 : (concat_22877 == 32'h0000_000a ? ____fsm_vvadd_impl_state_27 : (concat_22877 == 32'h0000_000b ? ____fsm_vvadd_impl_state_28 : (concat_22877 == 32'h0000_000c ? ____fsm_vvadd_impl_state_29 : (concat_22877 == 32'h0000_000d ? ____fsm_vvadd_impl_state_30 : (concat_22877 == 32'h0000_000e ? ____fsm_vvadd_impl_state_31 : __fsm_vvadd_impl_state_30_select_v1_in_recv_before_loop)))))))))))))));
  assign p0_stage_done = p0_all_active_inputs_valid & (out_not_pred | out_rdy);
  assign v0_in_select = nor_22913 ? v0_in : 32'h0000_0000;
  assign sign_ext_22957 = {32{__fsm_vvadd_impl_in_state_15}};
  assign v0_in_recv_value = v0_in_select & {32{__fsm_vvadd_impl_in_state_0}};
  assign v0_in_recv_value__1 = v0_in_select & {32{__fsm_vvadd_impl_in_state_1}};
  assign v0_in_recv_value__2 = v0_in_select & {32{__fsm_vvadd_impl_in_state_2}};
  assign v0_in_recv_value__3 = v0_in_select & {32{__fsm_vvadd_impl_in_state_3}};
  assign v0_in_recv_value__4 = v0_in_select & {32{__fsm_vvadd_impl_in_state_4}};
  assign v0_in_recv_value__5 = v0_in_select & {32{__fsm_vvadd_impl_in_state_5}};
  assign v0_in_recv_value__6 = v0_in_select & {32{__fsm_vvadd_impl_in_state_6}};
  assign v0_in_recv_value__7 = v0_in_select & {32{__fsm_vvadd_impl_in_state_7}};
  assign v0_in_recv_value__8 = v0_in_select & {32{__fsm_vvadd_impl_in_state_8}};
  assign v0_in_recv_value__9 = v0_in_select & {32{__fsm_vvadd_impl_in_state_9}};
  assign v0_in_recv_value__10 = v0_in_select & {32{__fsm_vvadd_impl_in_state_10}};
  assign v0_in_recv_value__11 = v0_in_select & {32{__fsm_vvadd_impl_in_state_11}};
  assign v0_in_recv_value__12 = v0_in_select & {32{__fsm_vvadd_impl_in_state_12}};
  assign v0_in_recv_value__13 = v0_in_select & {32{__fsm_vvadd_impl_in_state_13}};
  assign v0_in_recv_value__14 = v0_in_select & {32{__fsm_vvadd_impl_in_state_14}};
  assign v0_in_recv_value__15 = v0_in_select & sign_ext_22957;
  assign v1_in_recv_value = v1_in_select & sign_ext_22957;
  assign v1_in_recv_value__1 = v1_in_select & {32{__fsm_vvadd_impl_in_state_16}};
  assign v1_in_recv_value__2 = v1_in_select & {32{__fsm_vvadd_impl_in_state_17}};
  assign v1_in_recv_value__3 = v1_in_select & {32{__fsm_vvadd_impl_in_state_18}};
  assign v1_in_recv_value__4 = v1_in_select & {32{__fsm_vvadd_impl_in_state_19}};
  assign v1_in_recv_value__5 = v1_in_select & {32{__fsm_vvadd_impl_in_state_20}};
  assign v1_in_recv_value__6 = v1_in_select & {32{__fsm_vvadd_impl_in_state_21}};
  assign v1_in_recv_value__7 = v1_in_select & {32{__fsm_vvadd_impl_in_state_22}};
  assign v1_in_recv_value__8 = v1_in_select & {32{__fsm_vvadd_impl_in_state_23}};
  assign v1_in_recv_value__9 = v1_in_select & {32{__fsm_vvadd_impl_in_state_24}};
  assign v1_in_recv_value__10 = v1_in_select & {32{__fsm_vvadd_impl_in_state_25}};
  assign v1_in_recv_value__11 = v1_in_select & {32{__fsm_vvadd_impl_in_state_26}};
  assign v1_in_recv_value__12 = v1_in_select & {32{__fsm_vvadd_impl_in_state_27}};
  assign v1_in_recv_value__13 = v1_in_select & {32{__fsm_vvadd_impl_in_state_28}};
  assign v1_in_recv_value__14 = v1_in_select & {32{__fsm_vvadd_impl_in_state_29}};
  assign concat_23037 = {and_22972, __fsm_vvadd_impl_in_state_31, __fsm_vvadd_impl_in_state_32, __fsm_vvadd_impl_in_state_33, __fsm_vvadd_impl_in_state_34, __fsm_vvadd_impl_in_state_35, __fsm_vvadd_impl_in_state_36, __fsm_vvadd_impl_in_state_37, __fsm_vvadd_impl_in_state_38, __fsm_vvadd_impl_in_state_39, __fsm_vvadd_impl_in_state_40, __fsm_vvadd_impl_in_state_41, __fsm_vvadd_impl_in_state_42, __fsm_vvadd_impl_in_state_43, __fsm_vvadd_impl_in_state_44, __fsm_vvadd_impl_in_final_state};
  assign out_send_value__15 = ____for_1_c[4'hf];
  assign out_send_value__14 = ____for_1_c[4'he];
  assign out_send_value__13 = ____for_1_c[4'hd];
  assign out_send_value__12 = ____for_1_c[4'hc];
  assign out_send_value__11 = ____for_1_c[4'hb];
  assign out_send_value__10 = ____for_1_c[4'ha];
  assign out_send_value__9 = ____for_1_c[4'h9];
  assign out_send_value__8 = ____for_1_c[4'h8];
  assign out_send_value__7 = ____for_1_c[4'h7];
  assign out_send_value__6 = ____for_1_c[4'h6];
  assign out_send_value__5 = ____for_1_c[4'h5];
  assign out_send_value__4 = ____for_1_c[4'h4];
  assign out_send_value__3 = ____for_1_c[4'h3];
  assign out_send_value__2 = ____for_1_c[4'h2];
  assign out_send_value__1 = ____for_1_c[4'h1];
  assign out_send_value = array_update_22987[4'h0];
  assign ____fsm_vvadd_impl_state_0__at_most_one_next_value = nor_22917 == one_hot_22988[1] & and_22918 == one_hot_22988[0];
  assign concat_23234 = {nor_22917 & p0_stage_done, and_22918 & p0_stage_done};
  assign __fsm_vvadd_impl_state_plus_one = ____fsm_vvadd_impl_state_0 + __fsm_vvadd_impl_state_1_index;
  assign __fsm_vvadd_impl_state_0_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value : ____fsm_vvadd_impl_state_1;
  assign __fsm_vvadd_impl_state_1_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__1 : ____fsm_vvadd_impl_state_2;
  assign __fsm_vvadd_impl_state_2_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__2 : ____fsm_vvadd_impl_state_3;
  assign __fsm_vvadd_impl_state_3_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__3 : ____fsm_vvadd_impl_state_4;
  assign __fsm_vvadd_impl_state_4_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__4 : ____fsm_vvadd_impl_state_5;
  assign __fsm_vvadd_impl_state_5_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__5 : ____fsm_vvadd_impl_state_6;
  assign __fsm_vvadd_impl_state_6_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__6 : ____fsm_vvadd_impl_state_7;
  assign __fsm_vvadd_impl_state_7_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__7 : ____fsm_vvadd_impl_state_8;
  assign __fsm_vvadd_impl_state_8_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__8 : ____fsm_vvadd_impl_state_9;
  assign __fsm_vvadd_impl_state_9_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__9 : ____fsm_vvadd_impl_state_10;
  assign __fsm_vvadd_impl_state_10_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__10 : ____fsm_vvadd_impl_state_11;
  assign __fsm_vvadd_impl_state_11_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__11 : ____fsm_vvadd_impl_state_12;
  assign __fsm_vvadd_impl_state_12_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__12 : ____fsm_vvadd_impl_state_13;
  assign __fsm_vvadd_impl_state_13_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__13 : ____fsm_vvadd_impl_state_14;
  assign __fsm_vvadd_impl_state_14_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__14 : ____fsm_vvadd_impl_state_15;
  assign __fsm_vvadd_impl_state_15_select_v0_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v0_in_recv_value__15 : ____fsm_vvadd_impl_state_16;
  assign __fsm_vvadd_impl_state_15_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value : ____fsm_vvadd_impl_state_17;
  assign __fsm_vvadd_impl_state_16_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__1 : ____fsm_vvadd_impl_state_18;
  assign __fsm_vvadd_impl_state_17_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__2 : ____fsm_vvadd_impl_state_19;
  assign __fsm_vvadd_impl_state_18_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__3 : ____fsm_vvadd_impl_state_20;
  assign __fsm_vvadd_impl_state_19_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__4 : ____fsm_vvadd_impl_state_21;
  assign __fsm_vvadd_impl_state_20_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__5 : ____fsm_vvadd_impl_state_22;
  assign __fsm_vvadd_impl_state_21_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__6 : ____fsm_vvadd_impl_state_23;
  assign __fsm_vvadd_impl_state_22_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__7 : ____fsm_vvadd_impl_state_24;
  assign __fsm_vvadd_impl_state_23_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__8 : ____fsm_vvadd_impl_state_25;
  assign __fsm_vvadd_impl_state_24_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__9 : ____fsm_vvadd_impl_state_26;
  assign __fsm_vvadd_impl_state_25_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__10 : ____fsm_vvadd_impl_state_27;
  assign __fsm_vvadd_impl_state_26_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__11 : ____fsm_vvadd_impl_state_28;
  assign __fsm_vvadd_impl_state_27_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__12 : ____fsm_vvadd_impl_state_29;
  assign __fsm_vvadd_impl_state_28_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__13 : ____fsm_vvadd_impl_state_30;
  assign __fsm_vvadd_impl_state_29_select_v1_in_recv_before_loop = ____fsm_vvadd_impl_exited_last_activation ? v1_in_recv_value__14 : ____fsm_vvadd_impl_state_31;
  assign __for_1_guarded_update_state_elements = ~(~__fsm_vvadd_impl_in_state_30 | and_22811[4]);
  assign or_23326 = ~p0_stage_done | ____fsm_vvadd_impl_state_0__at_most_one_next_value | rst;
  assign one_hot_sel_23235 = __fsm_vvadd_impl_state_0_index & {6{concat_23234[0]}} | __fsm_vvadd_impl_state_plus_one & {6{concat_23234[1]}};
  assign and_23283 = (nor_22917 | and_22918) & p0_stage_done;
  assign sel_23095 = ____fsm_vvadd_impl_state_0 == 6'h00 ? __fsm_vvadd_impl_state_0_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h01 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h02 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h03 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h04 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h05 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h06 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h07 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h08 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h09 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h0a ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h0b ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h0c ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h0d ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h0e ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_1 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_1 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23096 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? __fsm_vvadd_impl_state_1_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h02 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h03 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h04 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h05 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h06 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h07 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h08 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h09 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h0a ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h0b ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h0c ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h0d ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h0e ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_2 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_2 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23097 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? __fsm_vvadd_impl_state_2_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h03 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h04 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h05 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h06 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h07 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h08 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h09 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h0a ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h0b ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h0c ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h0d ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h0e ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_3 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_3 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23098 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? __fsm_vvadd_impl_state_3_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h04 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h05 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h06 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h07 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h08 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h09 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h0a ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h0b ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h0c ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h0d ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h0e ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_4 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_4 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23099 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? __fsm_vvadd_impl_state_4_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h05 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h06 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h07 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h08 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h09 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h0a ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h0b ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h0c ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h0d ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h0e ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_5 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_5 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23100 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? __fsm_vvadd_impl_state_5_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h06 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h07 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h08 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h09 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h0a ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h0b ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h0c ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h0d ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h0e ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_6 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_6 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23101 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? __fsm_vvadd_impl_state_6_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h07 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h08 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h09 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h0a ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h0b ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h0c ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h0d ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h0e ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_7 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_7 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23102 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? __fsm_vvadd_impl_state_7_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h08 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h09 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h0a ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h0b ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h0c ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h0d ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h0e ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_8 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_8 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23103 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? __fsm_vvadd_impl_state_8_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h09 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h0a ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h0b ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h0c ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h0d ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h0e ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_9 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_9 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23104 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? __fsm_vvadd_impl_state_9_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h0a ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h0b ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h0c ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h0d ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h0e ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_10 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_10 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23105 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? __fsm_vvadd_impl_state_10_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h0b ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h0c ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h0d ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h0e ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_11 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_11 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23106 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? __fsm_vvadd_impl_state_11_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h0c ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h0d ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h0e ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_12 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_12 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23107 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? __fsm_vvadd_impl_state_12_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h0d ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h0e ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_13 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_13 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23108 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? __fsm_vvadd_impl_state_13_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h0e ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_14 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_14 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23109 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? __fsm_vvadd_impl_state_14_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h0f ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_15 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_15 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23110 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? __fsm_vvadd_impl_state_15_select_v0_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_16 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_16 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23111 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? __fsm_vvadd_impl_state_15_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h10 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_17 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_17 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23112 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? __fsm_vvadd_impl_state_16_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h11 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_18 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_18 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23113 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h11 ? __fsm_vvadd_impl_state_17_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h12 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_19 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_19 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23114 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h11 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h12 ? __fsm_vvadd_impl_state_18_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h13 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_20 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_20 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23115 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h11 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h12 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h13 ? __fsm_vvadd_impl_state_19_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h14 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_21 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_21 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23116 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h11 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h12 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h13 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h14 ? __fsm_vvadd_impl_state_20_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h15 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_22 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_22 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23117 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h11 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h12 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h13 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h14 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h15 ? __fsm_vvadd_impl_state_21_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h16 ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_23 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_23 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23118 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h11 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h12 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h13 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h14 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h15 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h16 ? __fsm_vvadd_impl_state_22_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h17 ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_24 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_24 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23119 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h11 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h12 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h13 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h14 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h15 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h16 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h17 ? __fsm_vvadd_impl_state_23_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h18 ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_25 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_25 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23120 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h11 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h12 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h13 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h14 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h15 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h16 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h17 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h18 ? __fsm_vvadd_impl_state_24_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h19 ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_26 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_26 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23121 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h11 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h12 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h13 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h14 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h15 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h16 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h17 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h18 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h19 ? __fsm_vvadd_impl_state_25_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h1a ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_27 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_27 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23122 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h11 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h12 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h13 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h14 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h15 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h16 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h17 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h18 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h19 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1a ? __fsm_vvadd_impl_state_26_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h1b ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_28 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_28 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23123 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h11 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h12 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h13 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h14 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h15 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h16 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h17 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h18 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h19 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1b ? __fsm_vvadd_impl_state_27_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h1c ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_29 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_29 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23124 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h11 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h12 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h13 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h14 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h15 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h16 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h17 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h18 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h19 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1c ? __fsm_vvadd_impl_state_28_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h1d ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_30 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_30 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23125 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h11 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h12 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h13 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h14 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h15 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h16 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h17 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h18 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h19 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1d ? __fsm_vvadd_impl_state_29_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h1e ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_31 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_31 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign sel_23126 = ____fsm_vvadd_impl_state_0 == 6'h00 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h01 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h02 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h03 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h04 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h05 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h06 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h07 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h08 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h09 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0e ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h0f ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h10 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h11 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h12 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h13 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h14 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h15 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h16 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h17 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h18 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h19 ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1a ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1b ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1c ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1d ? 32'h0000_0000 : (____fsm_vvadd_impl_state_0 == 6'h1e ? __fsm_vvadd_impl_state_30_select_v1_in_recv_before_loop : (____fsm_vvadd_impl_state_0 == 6'h1f ? ____fsm_vvadd_impl_state_32 : (____fsm_vvadd_impl_state_0 == 6'h20 ? ____fsm_vvadd_impl_state_32 : (____fsm_vvadd_impl_state_0 == 6'h21 ? ____fsm_vvadd_impl_state_32 : (____fsm_vvadd_impl_state_0 == 6'h22 ? ____fsm_vvadd_impl_state_32 : (____fsm_vvadd_impl_state_0 == 6'h23 ? ____fsm_vvadd_impl_state_32 : (____fsm_vvadd_impl_state_0 == 6'h24 ? ____fsm_vvadd_impl_state_32 : (____fsm_vvadd_impl_state_0 == 6'h25 ? ____fsm_vvadd_impl_state_32 : (____fsm_vvadd_impl_state_0 == 6'h26 ? ____fsm_vvadd_impl_state_32 : (____fsm_vvadd_impl_state_0 == 6'h27 ? ____fsm_vvadd_impl_state_32 : (____fsm_vvadd_impl_state_0 == 6'h28 ? ____fsm_vvadd_impl_state_32 : (____fsm_vvadd_impl_state_0 == 6'h29 ? ____fsm_vvadd_impl_state_32 : (____fsm_vvadd_impl_state_0 == 6'h2a ? ____fsm_vvadd_impl_state_32 : (____fsm_vvadd_impl_state_0 == 6'h2b ? ____fsm_vvadd_impl_state_32 : (____fsm_vvadd_impl_state_0 == 6'h2c ? ____fsm_vvadd_impl_state_32 : (____fsm_vvadd_impl_state_0 == 6'h2d ? ____fsm_vvadd_impl_state_32 : 32'h0000_0000)))))))))))))))))))))))))))))))))))))))))))));
  assign and_23317 = __fsm_vvadd_impl_in_state_30 & p0_stage_done;
  assign and_23319 = __for_1_guarded_update_state_elements & p0_stage_done;
  assign unexpand_for___for_1_i_next__1_case_1 = add_22847[4:0];
  always_ff @ (posedge clk) begin
    if (rst) begin
      ____for_1__last_iter_broke <= 1'h1;
      ____fsm_vvadd_impl_state_0 <= 6'h00;
      ____for_1_i <= 5'h00;
      ____fsm_vvadd_impl_exited_last_activation <= 1'h1;
      ____fsm_vvadd_impl_state_32 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_1 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_2 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_3 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_4 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_5 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_6 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_7 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_8 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_9 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_10 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_11 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_12 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_13 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_14 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_15 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_16 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_17 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_18 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_19 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_20 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_21 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_22 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_23 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_24 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_25 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_26 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_27 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_28 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_29 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_30 <= 32'h0000_0000;
      ____fsm_vvadd_impl_state_31 <= 32'h0000_0000;
      ____for_1_c <= ____for_1_c_init;
    end else begin
      ____for_1__last_iter_broke <= and_23317 ? __for_1_do_break_from_func : ____for_1__last_iter_broke;
      ____fsm_vvadd_impl_state_0 <= and_23283 ? one_hot_sel_23235 : ____fsm_vvadd_impl_state_0;
      ____for_1_i <= and_23319 ? unexpand_for___for_1_i_next__1_case_1 : ____for_1_i;
      ____fsm_vvadd_impl_exited_last_activation <= p0_stage_done ? __fsm_vvadd_impl_go_to_next_state_in_state : ____fsm_vvadd_impl_exited_last_activation;
      ____fsm_vvadd_impl_state_32 <= p0_stage_done ? sel_23126 : ____fsm_vvadd_impl_state_32;
      ____fsm_vvadd_impl_state_1 <= p0_stage_done ? sel_23095 : ____fsm_vvadd_impl_state_1;
      ____fsm_vvadd_impl_state_2 <= p0_stage_done ? sel_23096 : ____fsm_vvadd_impl_state_2;
      ____fsm_vvadd_impl_state_3 <= p0_stage_done ? sel_23097 : ____fsm_vvadd_impl_state_3;
      ____fsm_vvadd_impl_state_4 <= p0_stage_done ? sel_23098 : ____fsm_vvadd_impl_state_4;
      ____fsm_vvadd_impl_state_5 <= p0_stage_done ? sel_23099 : ____fsm_vvadd_impl_state_5;
      ____fsm_vvadd_impl_state_6 <= p0_stage_done ? sel_23100 : ____fsm_vvadd_impl_state_6;
      ____fsm_vvadd_impl_state_7 <= p0_stage_done ? sel_23101 : ____fsm_vvadd_impl_state_7;
      ____fsm_vvadd_impl_state_8 <= p0_stage_done ? sel_23102 : ____fsm_vvadd_impl_state_8;
      ____fsm_vvadd_impl_state_9 <= p0_stage_done ? sel_23103 : ____fsm_vvadd_impl_state_9;
      ____fsm_vvadd_impl_state_10 <= p0_stage_done ? sel_23104 : ____fsm_vvadd_impl_state_10;
      ____fsm_vvadd_impl_state_11 <= p0_stage_done ? sel_23105 : ____fsm_vvadd_impl_state_11;
      ____fsm_vvadd_impl_state_12 <= p0_stage_done ? sel_23106 : ____fsm_vvadd_impl_state_12;
      ____fsm_vvadd_impl_state_13 <= p0_stage_done ? sel_23107 : ____fsm_vvadd_impl_state_13;
      ____fsm_vvadd_impl_state_14 <= p0_stage_done ? sel_23108 : ____fsm_vvadd_impl_state_14;
      ____fsm_vvadd_impl_state_15 <= p0_stage_done ? sel_23109 : ____fsm_vvadd_impl_state_15;
      ____fsm_vvadd_impl_state_16 <= p0_stage_done ? sel_23110 : ____fsm_vvadd_impl_state_16;
      ____fsm_vvadd_impl_state_17 <= p0_stage_done ? sel_23111 : ____fsm_vvadd_impl_state_17;
      ____fsm_vvadd_impl_state_18 <= p0_stage_done ? sel_23112 : ____fsm_vvadd_impl_state_18;
      ____fsm_vvadd_impl_state_19 <= p0_stage_done ? sel_23113 : ____fsm_vvadd_impl_state_19;
      ____fsm_vvadd_impl_state_20 <= p0_stage_done ? sel_23114 : ____fsm_vvadd_impl_state_20;
      ____fsm_vvadd_impl_state_21 <= p0_stage_done ? sel_23115 : ____fsm_vvadd_impl_state_21;
      ____fsm_vvadd_impl_state_22 <= p0_stage_done ? sel_23116 : ____fsm_vvadd_impl_state_22;
      ____fsm_vvadd_impl_state_23 <= p0_stage_done ? sel_23117 : ____fsm_vvadd_impl_state_23;
      ____fsm_vvadd_impl_state_24 <= p0_stage_done ? sel_23118 : ____fsm_vvadd_impl_state_24;
      ____fsm_vvadd_impl_state_25 <= p0_stage_done ? sel_23119 : ____fsm_vvadd_impl_state_25;
      ____fsm_vvadd_impl_state_26 <= p0_stage_done ? sel_23120 : ____fsm_vvadd_impl_state_26;
      ____fsm_vvadd_impl_state_27 <= p0_stage_done ? sel_23121 : ____fsm_vvadd_impl_state_27;
      ____fsm_vvadd_impl_state_28 <= p0_stage_done ? sel_23122 : ____fsm_vvadd_impl_state_28;
      ____fsm_vvadd_impl_state_29 <= p0_stage_done ? sel_23123 : ____fsm_vvadd_impl_state_29;
      ____fsm_vvadd_impl_state_30 <= p0_stage_done ? sel_23124 : ____fsm_vvadd_impl_state_30;
      ____fsm_vvadd_impl_state_31 <= p0_stage_done ? sel_23125 : ____fsm_vvadd_impl_state_31;
      ____for_1_c <= and_23319 ? array_update_22987 : ____for_1_c;
    end
  end
  assign out = out_send_value__15 & {32{concat_23037[0]}} | out_send_value__14 & {32{concat_23037[1]}} | out_send_value__13 & {32{concat_23037[2]}} | out_send_value__12 & {32{concat_23037[3]}} | out_send_value__11 & {32{concat_23037[4]}} | out_send_value__10 & {32{concat_23037[5]}} | out_send_value__9 & {32{concat_23037[6]}} | out_send_value__8 & {32{concat_23037[7]}} | out_send_value__7 & {32{concat_23037[8]}} | out_send_value__6 & {32{concat_23037[9]}} | out_send_value__5 & {32{concat_23037[10]}} | out_send_value__4 & {32{concat_23037[11]}} | out_send_value__3 & {32{concat_23037[12]}} | out_send_value__2 & {32{concat_23037[13]}} | out_send_value__1 & {32{concat_23037[14]}} | out_send_value & {32{concat_23037[15]}};
  assign out_vld = p0_all_active_inputs_valid & or_23090;
  assign v0_in_rdy = p0_stage_done & nor_22913;
  assign v1_in_rdy = p0_stage_done & or_22846;
  for (genvar __i0 = 0; __i0 < 16; __i0 = __i0 + 1) begin : gen__array_update_22987_0
    assign array_update_22987[__i0] = concat_22877 == __i0 ? add_22939 : sel_22938[__i0];
  end
  `ifdef ASSERT_ON
  ____fsm_vvadd_impl_state_0__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_23326))) or_23326) else $fatal(0, "More than one next_value fired for state element: __fsm_vvadd_impl_state_0");
  `endif  // ASSERT_ON
endmodule
