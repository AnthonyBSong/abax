module mv_mem(
  input wire clk,
  input wire rst,
  input wire out_rdy,
  input wire v0__read_req_rdy,
  input wire [31:0] v0__read_resp,
  input wire v0__read_resp_vld,
  input wire v0__write_completion_vld,
  input wire v0__write_req_rdy,
  input wire [31:0] v0_in,
  input wire v0_in_vld,
  input wire v1__read_req_rdy,
  input wire [31:0] v1__read_resp,
  input wire v1__read_resp_vld,
  input wire v1__write_completion_vld,
  input wire v1__write_req_rdy,
  input wire [31:0] v1_in,
  input wire v1_in_vld,
  input wire [31:0] y_rd_data,
  output wire [31:0] out,
  output wire out_vld,
  output wire [3:0] v0__read_req,
  output wire v0__read_req_vld,
  output wire v0__read_resp_rdy,
  output wire v0__write_completion_rdy,
  output wire [35:0] v0__write_req,
  output wire v0__write_req_vld,
  output wire v0_in_rdy,
  output wire [1:0] v1__read_req,
  output wire v1__read_req_vld,
  output wire v1__read_resp_rdy,
  output wire v1__write_completion_rdy,
  output wire [33:0] v1__write_req,
  output wire v1__write_req_vld,
  output wire v1_in_rdy,
  output wire [1:0] y_rd_addr,
  output wire y_rd_en,
  output wire [1:0] y_wr_addr,
  output wire [31:0] y_wr_data,
  output wire y_wr_en
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] smul32b_32b_x_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    reg signed [31:0] signed_lhs;
    reg signed [31:0] signed_rhs;
    reg signed [31:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul32b_32b_x_32b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  wire [31:0] literal_5840 = 32'h0000_0000;
  wire [31:0] literal_5756 = 32'h0000_0000;
  wire [31:0] literal_5760 = 32'h0000_0000;
  wire [1:0] literal_5421[4];
  assign literal_5421 = '{2'h1, 2'h2, 2'h3, 2'h0};
  reg ____for_4__last_iter_broke;
  reg ____for_2__last_iter_broke;
  reg ____for_3__last_iter_broke;
  reg ____for_5__last_iter_broke;
  reg ____for_1__last_iter_broke;
  reg [5:0] ____for_4_j;
  reg [2:0] ____for_2__i;
  reg [5:0] ____for_3_i;
  reg [2:0] ____for_5__i;
  reg [4:0] ____for_1__i;
  reg [2:0] ____fsm_mv_impl_state;
  reg [1:0] __this;
  reg ____fsm___for_3_loop_state;
  reg ____fsm___for_4_loop_state_0;
  reg p0_____fsm___for_4_loop_state_0__1;
  reg p0___fsm_mv_impl_in_state_1;
  reg p0___for_2_loop_contents_condition;
  reg p0_ctx_5__full_condition_ctx_6__ful_output;
  reg p0___fsm___for_4_loop_in_state_0;
  reg p0___fsm___for_4_loop_returns_this_activation_vars;
  reg p0___for_5_loop_contents_condition;
  reg p0___fsm_mv_impl_in_state_2;
  reg p0___fsm_mv_impl_in_state_3;
  reg p0___fsm_mv_impl_in_state_4;
  reg p0_and_5554;
  reg p0___for_1_loop_contents_condition;
  reg p0_nor_5558;
  reg p0_not_5663;
  reg [1:0] p0_tuple_5586_index0;
  reg p0_nand_5664;
  reg p0_nand_5665;
  reg p0_and_5582;
  reg p0_and_5583;
  reg [31:0] ____fsm___for_4_loop_state_1;
  reg [31:0] ____fsm___for_4_loop_state_2;
  reg p1_____fsm___for_4_loop_state_0__1;
  reg p1___fsm_mv_impl_in_state_1;
  reg p1_ctx_5__full_condition_ctx_6__ful_output;
  reg [31:0] p1_smul_5746;
  reg p1___fsm___for_4_loop_in_state_0;
  reg p1___fsm___for_4_loop_returns_this_activation_vars;
  reg p1___for_5_loop_contents_condition;
  reg p1___fsm_mv_impl_in_state_2;
  reg p1___fsm_mv_impl_in_state_3;
  reg p1___fsm_mv_impl_in_state_4;
  reg p1_and_5554;
  reg p1_nor_5558;
  reg p1_not_5663;
  reg p1_not_5767;
  reg p1_or_5748;
  reg p1_nand_5664;
  reg p1_nand_5665;
  reg p1_and_5582;
  reg p1_and_5583;
  reg [31:0] ____fsm___for_4_loop_state_3;
  reg p2___fsm___for_4_loop_returns_this_activation_vars;
  reg p2_nor_5558;
  reg p2_and_5834;
  reg p2_and_5818;
  reg p2_and_5817;
  reg p2_and_5816;
  reg p2_not_5663;
  reg p2_or_5838;
  reg p2_nand_5665;
  reg p2_nand_5851;
  reg p2_nand_5852;
  reg p2_nand_5853;
  reg p2_nand_5854;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg __v1__write_req_has_been_sent_reg;
  reg __v0__read_req_has_been_sent_reg;
  reg __v1__read_req_has_been_sent_reg;
  reg __v0__write_req_has_been_sent_reg;
  reg __y__read_req_has_been_sent_reg;
  reg __y__write_req_has_been_sent_reg;
  reg __out_has_been_sent_reg;
  reg __y_rd_en__1_delay_reg;
  reg [31:0] __y_ram_zero_latency0_skid_reg;
  reg __y_ram_zero_latency0_valid_skid_reg;
  wire __fsm___for_4_loop_default_next_state;
  wire [5:0] and_5505;
  wire [2:0] and_5510;
  wire [5:0] and_5511;
  wire [2:0] __fsm_mv_impl_state_5_index;
  wire [2:0] and_5515;
  wire [4:0] and_5516;
  wire [6:0] add_5519;
  wire __fsm_mv_impl_in_state_5;
  wire ctx_5__full_condition_ctx_6__ful_output;
  wire [3:0] add_5527;
  wire [6:0] add_5528;
  wire [1:0] __fsm___for_3_loop_initial_state_index;
  wire __fsm___for_4_loop_go_to_next_state;
  wire [3:0] add_5532;
  wire [5:0] add_5534;
  wire __for_4_do_break_from_func;
  wire __fsm___for_4_loop_returns_this_activation_vars;
  wire __for_2_do_break_from_func;
  wire __for_3_do_break_from_func;
  wire __for_4_do_break_with_fsm;
  wire __for_5_do_break_from_func;
  wire [2:0] __fsm_mv_impl_state_0_index;
  wire __for_1_do_break_from_func;
  wire ctx_5__full_condition_continuati_output;
  wire __for_3_not_enter_condition;
  wire __for_3_do_break_with_fsm;
  wire ctx_6__full_condition_continuati_output;
  wire [2:0] __fsm_mv_impl_state_1_index;
  wire __fsm_mv_impl_in_state_0;
  wire __for_1_not_exit_state_condition;
  wire __for_2_not_exit_state_condition;
  wire __for_4_enter_condition;
  wire __for_3_not_exit_state_condition;
  wire __for_5_not_exit_state_condition;
  wire not_5904;
  wire or_5748;
  wire __fsm_mv_impl_in_state_1;
  wire __fsm___for_4_loop_in_state_0;
  wire __fsm_mv_impl_go_to_next_state_in_state;
  wire [2:0] __fsm_mv_impl_state_6_index;
  wire or_6245;
  wire p2_all_active_outputs_ready;
  wire y__read_req_not_pred;
  wire y_ram_zero_latency0_from_skid_rdy;
  wire __for_2_loop_contents_condition;
  wire __for_1_loop_contents_condition;
  wire and_5554;
  wire __fsm_mv_impl_in_state_6;
  wire p2_stage_done;
  wire p2_not_valid;
  wire p1_all_active_inputs_valid;
  wire or_6251;
  wire v0__read_req_not_pred;
  wire nor_5593;
  wire __fsm_mv_impl_returns_this_activation_vars;
  wire nor_5558;
  wire p1_enable;
  wire p1_stage_done;
  wire [1:0] ____fsm_mv_impl_state__next_value_predicates;
  wire [1:0] ____fsm___for_3_loop_state__next_value_predicates;
  wire [1:0] ____fsm___for_4_loop_state_0__next_value_predicates;
  wire p1_data_enable;
  wire p1_not_valid;
  wire p0_all_active_inputs_valid;
  wire p0_all_active_outputs_ready;
  wire [31:0] y_ram_zero_latency0_select;
  wire [2:0] one_hot_5607;
  wire [2:0] one_hot_5608;
  wire [2:0] one_hot_5609;
  wire p0_enable;
  wire p0_stage_done;
  wire and_5834;
  wire and_5818;
  wire and_5817;
  wire and_5816;
  wire [1:0] y_read_addr;
  wire p0_data_enable;
  wire __v1__write_req_vld_buf;
  wire __v1__write_req_not_has_been_sent;
  wire __v0__read_req_vld_buf;
  wire __v0__read_req_not_has_been_sent;
  wire __v1__read_req_not_has_been_sent;
  wire __v0__write_req_vld_buf;
  wire __v0__write_req_not_has_been_sent;
  wire __y__read_req_vld_buf;
  wire __y__read_req_not_has_been_sent;
  wire or_5838;
  wire __out_vld_buf;
  wire __out_not_has_been_sent;
  wire and_6109;
  wire [31:0] y_write_value__5;
  wire [31:0] y__read_resp_select;
  wire [1:0] add_5588;
  wire [1:0] v1_read_addr;
  wire __for_5_loop_contents_condition;
  wire and_6033;
  wire and_6034;
  wire and_6082;
  wire and_6083;
  wire and_6089;
  wire and_6090;
  wire __v1__write_req_valid_and_not_has_been_sent;
  wire __v0__read_req_valid_and_not_has_been_sent;
  wire __v1__read_req_valid_and_not_has_been_sent;
  wire __v0__write_req_valid_and_not_has_been_sent;
  wire y_rd_en__1;
  wire __y__write_req_vld_buf;
  wire __y__write_req_not_has_been_sent;
  wire __out_valid_and_not_has_been_sent;
  wire y_ram_zero_latency0_to_is_not_rdy;
  wire [31:0] tuple_index_5845;
  wire [3:0] v0_read_addr;
  wire [3:0] v0_write_addr;
  wire [31:0] v0_in_select;
  wire [1:0] v1_write_addr;
  wire [31:0] v1_in_select;
  wire ____fsm_mv_impl_state__at_most_one_next_value;
  wire ____fsm___for_3_loop_state__at_most_one_next_value;
  wire ____fsm___for_4_loop_state_0__at_most_one_next_value;
  wire [2:0] __fsm_mv_impl_state_2_index;
  wire [2:0] __fsm_mv_impl_state_3_index;
  wire [2:0] __fsm_mv_impl_state_4_index;
  wire [1:0] concat_5565;
  wire [1:0] y_read_addr__1;
  wire or_5572;
  wire [1:0] concat_6036;
  wire [2:0] __fsm_mv_impl_state_plus_one;
  wire [31:0] v0__read_resp_select;
  wire [31:0] v1__read_resp_select;
  wire continuation_1_ctx_3__full_condi_output;
  wire __for_1_initial_loop_cond;
  wire __for_2_guarded_update_state_elements;
  wire __for_3_initial_loop_cond;
  wire __for_4_initial_loop_cond;
  wire __for_5_guarded_update_state_elements;
  wire [1:0] concat_6085;
  wire [1:0] concat_6092;
  wire __v1__write_req_valid_and_all_active_outputs_ready;
  wire __v1__write_req_valid_and_ready_txfr;
  wire __v0__read_req_valid_and_all_active_outputs_ready;
  wire __v0__read_req_valid_and_ready_txfr;
  wire __v1__read_req_valid_and_ready_txfr;
  wire __v0__write_req_valid_and_all_active_outputs_ready;
  wire __v0__write_req_valid_and_ready_txfr;
  wire __y__read_req_valid_and_all_active_outputs_ready;
  wire __y__read_req_valid_and_ready_txfr;
  wire __y__write_req_valid_and_all_active_outputs_ready;
  wire y_wr_en__1;
  wire __out_valid_and_all_active_outputs_ready;
  wire __out_valid_and_ready_txfr;
  wire y_ram_zero_latency0_skid_data_load_en;
  wire y_ram_zero_latency0_skid_valid_set_zero;
  wire [1:0] tuple_5733;
  wire [33:0] tuple_5837;
  wire [31:0] y_read_response__1;
  wire and_6103;
  wire and_6105;
  wire and_6108;
  wire or_6240;
  wire or_6242;
  wire or_6244;
  wire p3_enable;
  wire p2_enable;
  wire nand_5851;
  wire nand_5852;
  wire nand_5853;
  wire nand_5854;
  wire [31:0] smul_5746;
  wire __fsm_mv_impl_in_state_2;
  wire __fsm_mv_impl_in_state_3;
  wire __fsm_mv_impl_in_state_4;
  wire not_5663;
  wire [1:0] one_hot_sel_5580;
  wire nand_5664;
  wire nand_5665;
  wire and_5582;
  wire and_5583;
  wire [2:0] one_hot_sel_6037;
  wire or_6038;
  wire [31:0] v0_read_response;
  wire and_6052;
  wire [31:0] v1_read_response;
  wire [31:0] y_read_response;
  wire and_6058;
  wire and_6061;
  wire [1:0] unexpand_for_this_next__1_case_1;
  wire [4:0] unexpand_for___for_1__i_next__1_case_1;
  wire and_6261;
  wire [2:0] unexpand_for___for_2__i_next__1_case_1;
  wire and_6070;
  wire [5:0] unexpand_for___for_3_i_next__1_case_1;
  wire and_6262;
  wire [5:0] unexpand_for___for_4_j_next__1_case_1;
  wire and_6263;
  wire [2:0] unexpand_for___for_5__i_next__1_case_1;
  wire and_6079;
  wire one_hot_sel_6086;
  wire or_6087;
  wire one_hot_sel_6093;
  wire or_6094;
  wire __v1__write_req_not_stage_load;
  wire __v1__write_req_has_been_sent_reg_load_en;
  wire __v0__read_req_not_stage_load;
  wire __v0__read_req_has_been_sent_reg_load_en;
  wire __v1__read_req_has_been_sent_reg_load_en;
  wire __v0__write_req_not_stage_load;
  wire __v0__write_req_has_been_sent_reg_load_en;
  wire __y__read_req_not_stage_load;
  wire __y__read_req_has_been_sent_reg_load_en;
  wire __y__write_req_not_stage_load;
  wire __y__write_req_has_been_sent_reg_load_en;
  wire __out_not_stage_load;
  wire __out_has_been_sent_reg_load_en;
  wire y_ram_zero_latency0_skid_valid_load_en;
  assign __fsm___for_4_loop_default_next_state = 1'h0;
  assign and_5505 = {6{~____for_4__last_iter_broke}} & ____for_4_j;
  assign and_5510 = {3{~____for_2__last_iter_broke}} & ____for_2__i;
  assign and_5511 = {6{~____for_3__last_iter_broke}} & ____for_3_i;
  assign __fsm_mv_impl_state_5_index = 3'h5;
  assign and_5515 = {3{~____for_5__last_iter_broke}} & ____for_5__i;
  assign and_5516 = {5{~____for_1__last_iter_broke}} & ____for_1__i;
  assign add_5519 = {__fsm___for_4_loop_default_next_state, and_5505} + 7'h01;
  assign __fsm_mv_impl_in_state_5 = ____fsm_mv_impl_state == __fsm_mv_impl_state_5_index;
  assign ctx_5__full_condition_ctx_6__ful_output = __this == 2'h2;
  assign add_5527 = {__fsm___for_4_loop_default_next_state, and_5510} + 4'h1;
  assign add_5528 = {__fsm___for_4_loop_default_next_state, and_5511} + 7'h01;
  assign __fsm___for_3_loop_initial_state_index = 2'h0;
  assign __fsm___for_4_loop_go_to_next_state = __fsm_mv_impl_in_state_5 & ctx_5__full_condition_ctx_6__ful_output & ____fsm___for_3_loop_state;
  assign add_5532 = {__fsm___for_4_loop_default_next_state, and_5515} + 4'h1;
  assign add_5534 = {__fsm___for_4_loop_default_next_state, and_5516} + 6'h01;
  assign __for_4_do_break_from_func = add_5519[6:5] != __fsm___for_3_loop_initial_state_index;
  assign __fsm___for_4_loop_returns_this_activation_vars = __fsm___for_4_loop_go_to_next_state & ____fsm___for_4_loop_state_0;
  assign __for_2_do_break_from_func = add_5527[3:2] != __fsm___for_3_loop_initial_state_index;
  assign __for_3_do_break_from_func = add_5528[6:5] != __fsm___for_3_loop_initial_state_index;
  assign __for_4_do_break_with_fsm = __for_4_do_break_from_func & __fsm___for_4_loop_returns_this_activation_vars;
  assign __for_5_do_break_from_func = add_5532[3:2] != __fsm___for_3_loop_initial_state_index;
  assign __fsm_mv_impl_state_0_index = 3'h0;
  assign __for_1_do_break_from_func = add_5534[5:4] != __fsm___for_3_loop_initial_state_index;
  assign ctx_5__full_condition_continuati_output = __this == 2'h1;
  assign __for_3_not_enter_condition = ~ctx_5__full_condition_ctx_6__ful_output;
  assign __for_3_do_break_with_fsm = __for_3_do_break_from_func & __for_4_do_break_with_fsm;
  assign ctx_6__full_condition_continuati_output = __this == 2'h3;
  assign __fsm_mv_impl_state_1_index = 3'h1;
  assign __fsm_mv_impl_in_state_0 = ____fsm_mv_impl_state == __fsm_mv_impl_state_0_index;
  assign __for_1_not_exit_state_condition = __this[0] | __this[1] | __for_1_do_break_from_func;
  assign __for_2_not_exit_state_condition = ~(ctx_5__full_condition_continuati_output & ~__for_2_do_break_from_func);
  assign __for_4_enter_condition = 1'h1;
  assign __for_3_not_exit_state_condition = __for_3_not_enter_condition | __for_3_do_break_with_fsm;
  assign __for_5_not_exit_state_condition = ~(ctx_6__full_condition_continuati_output & ~__for_5_do_break_from_func);
  assign not_5904 = ~p0_and_5554;
  assign or_5748 = p0_and_5554 | p0___for_5_loop_contents_condition;
  assign __fsm_mv_impl_in_state_1 = ____fsm_mv_impl_state == __fsm_mv_impl_state_1_index;
  assign __fsm___for_4_loop_in_state_0 = ~____fsm___for_4_loop_state_0;
  assign __fsm_mv_impl_go_to_next_state_in_state = ____fsm_mv_impl_state == 3'h0 ? __for_1_not_exit_state_condition : (____fsm_mv_impl_state == 3'h1 ? __for_2_not_exit_state_condition : (____fsm_mv_impl_state == 3'h2 ? __for_4_enter_condition : (____fsm_mv_impl_state == 3'h3 ? __for_4_enter_condition : (____fsm_mv_impl_state == 3'h4 ? __for_4_enter_condition : (____fsm_mv_impl_state == 3'h5 ? __for_3_not_exit_state_condition : (____fsm_mv_impl_state == 3'h6 ? __for_5_not_exit_state_condition : __fsm___for_4_loop_default_next_state))))));
  assign __fsm_mv_impl_state_6_index = 3'h6;
  assign or_6245 = ~p1_or_5748 | __y_rd_en__1_delay_reg | __y_ram_zero_latency0_valid_skid_reg;
  assign p2_all_active_outputs_ready = ~p1___for_5_loop_contents_condition | out_rdy | __out_has_been_sent_reg;
  assign y__read_req_not_pred = ~or_5748;
  assign y_ram_zero_latency0_from_skid_rdy = ~__y_ram_zero_latency0_valid_skid_reg;
  assign __for_2_loop_contents_condition = __fsm_mv_impl_in_state_1 & ctx_5__full_condition_continuati_output;
  assign __for_1_loop_contents_condition = ~(~__fsm_mv_impl_in_state_0 | __this[0] | __this[1]);
  assign and_5554 = __fsm___for_4_loop_go_to_next_state & __fsm___for_4_loop_in_state_0;
  assign __fsm_mv_impl_in_state_6 = ____fsm_mv_impl_state == __fsm_mv_impl_state_6_index;
  assign p2_stage_done = p1_valid & or_6245 & p2_all_active_outputs_ready;
  assign p2_not_valid = ~p1_valid;
  assign p1_all_active_inputs_valid = (~p0___for_2_loop_contents_condition | v1__write_completion_vld) & (not_5904 | v0__read_resp_vld) & (not_5904 | v1__read_resp_vld) & (~p0___for_1_loop_contents_condition | v0__write_completion_vld);
  assign or_6251 = y__read_req_not_pred | y_ram_zero_latency0_from_skid_rdy | __y__read_req_has_been_sent_reg;
  assign v0__read_req_not_pred = ~and_5554;
  assign nor_5593 = ~(~__fsm_mv_impl_go_to_next_state_in_state | __fsm_mv_impl_in_state_6);
  assign __fsm_mv_impl_returns_this_activation_vars = __fsm_mv_impl_in_state_6 & __fsm_mv_impl_go_to_next_state_in_state;
  assign nor_5558 = ~(~__fsm_mv_impl_in_state_5 | __for_3_not_enter_condition | ____fsm___for_3_loop_state);
  assign p1_enable = p2_stage_done | p2_not_valid;
  assign p1_stage_done = p0_valid & p1_all_active_inputs_valid & or_6251;
  assign ____fsm_mv_impl_state__next_value_predicates = {nor_5593, __fsm_mv_impl_returns_this_activation_vars};
  assign ____fsm___for_3_loop_state__next_value_predicates = {nor_5558, __for_4_do_break_with_fsm};
  assign ____fsm___for_4_loop_state_0__next_value_predicates = {and_5554, __fsm___for_4_loop_returns_this_activation_vars};
  assign p1_data_enable = p1_enable & p1_stage_done;
  assign p1_not_valid = ~p0_valid;
  assign p0_all_active_inputs_valid = (~__for_2_loop_contents_condition | v1_in_vld) & (~__for_1_loop_contents_condition | v0_in_vld);
  assign p0_all_active_outputs_ready = (~__for_2_loop_contents_condition | v1__write_req_rdy | __v1__write_req_has_been_sent_reg) & (v0__read_req_not_pred | v0__read_req_rdy | __v0__read_req_has_been_sent_reg) & (v0__read_req_not_pred | v1__read_req_rdy | __v1__read_req_has_been_sent_reg) & (~__for_1_loop_contents_condition | v0__write_req_rdy | __v0__write_req_has_been_sent_reg);
  assign y_ram_zero_latency0_select = __y_ram_zero_latency0_valid_skid_reg ? __y_ram_zero_latency0_skid_reg : y_rd_data;
  assign one_hot_5607 = {____fsm_mv_impl_state__next_value_predicates[1:0] == 2'h0, ____fsm_mv_impl_state__next_value_predicates[1] && !____fsm_mv_impl_state__next_value_predicates[0], ____fsm_mv_impl_state__next_value_predicates[0]};
  assign one_hot_5608 = {____fsm___for_3_loop_state__next_value_predicates[1:0] == 2'h0, ____fsm___for_3_loop_state__next_value_predicates[1] && !____fsm___for_3_loop_state__next_value_predicates[0], ____fsm___for_3_loop_state__next_value_predicates[0]};
  assign one_hot_5609 = {____fsm___for_4_loop_state_0__next_value_predicates[1:0] == 2'h0, ____fsm___for_4_loop_state_0__next_value_predicates[1] && !____fsm___for_4_loop_state_0__next_value_predicates[0], ____fsm___for_4_loop_state_0__next_value_predicates[0]};
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign p0_stage_done = p0_all_active_inputs_valid & p0_all_active_outputs_ready;
  assign and_5834 = p1_ctx_5__full_condition_ctx_6__ful_output & p1___fsm_mv_impl_in_state_1;
  assign and_5818 = p1_ctx_5__full_condition_ctx_6__ful_output & p1___fsm_mv_impl_in_state_2;
  assign and_5817 = p1_ctx_5__full_condition_ctx_6__ful_output & p1___fsm_mv_impl_in_state_3;
  assign and_5816 = p1_ctx_5__full_condition_ctx_6__ful_output & p1___fsm_mv_impl_in_state_4;
  assign y_read_addr = and_5511[1:0];
  assign p0_data_enable = p0_enable & p0_stage_done;
  assign __v1__write_req_vld_buf = p0_all_active_inputs_valid & p0_enable & __for_2_loop_contents_condition;
  assign __v1__write_req_not_has_been_sent = ~__v1__write_req_has_been_sent_reg;
  assign __v0__read_req_vld_buf = p0_all_active_inputs_valid & p0_enable & and_5554;
  assign __v0__read_req_not_has_been_sent = ~__v0__read_req_has_been_sent_reg;
  assign __v1__read_req_not_has_been_sent = ~__v1__read_req_has_been_sent_reg;
  assign __v0__write_req_vld_buf = p0_all_active_inputs_valid & p0_enable & __for_1_loop_contents_condition;
  assign __v0__write_req_not_has_been_sent = ~__v0__write_req_has_been_sent_reg;
  assign __y__read_req_vld_buf = p1_all_active_inputs_valid & p0_valid & p1_enable & or_5748;
  assign __y__read_req_not_has_been_sent = ~__y__read_req_has_been_sent_reg;
  assign or_5838 = p1___fsm___for_4_loop_returns_this_activation_vars | p1_nor_5558 | and_5834 | and_5818 | and_5817 | and_5816;
  assign __out_vld_buf = or_6245 & p1_valid & p1___for_5_loop_contents_condition;
  assign __out_not_has_been_sent = ~__out_has_been_sent_reg;
  assign and_6109 = p2_stage_done & p1_or_5748;
  assign y_write_value__5 = ____fsm___for_4_loop_state_3 + p1_smul_5746;
  assign y__read_resp_select = p1_or_5748 ? {y_ram_zero_latency0_select} : literal_5840;
  assign add_5588 = y_read_addr + and_5505[3:2];
  assign v1_read_addr = and_5505[1:0];
  assign __for_5_loop_contents_condition = __fsm_mv_impl_in_state_6 & ctx_6__full_condition_continuati_output;
  assign and_6033 = nor_5593 & p0_data_enable;
  assign and_6034 = __fsm_mv_impl_returns_this_activation_vars & p0_data_enable;
  assign and_6082 = nor_5558 & p0_data_enable;
  assign and_6083 = __for_4_do_break_with_fsm & p0_data_enable;
  assign and_6089 = and_5554 & p0_data_enable;
  assign and_6090 = __fsm___for_4_loop_returns_this_activation_vars & p0_data_enable;
  assign __v1__write_req_valid_and_not_has_been_sent = __v1__write_req_vld_buf & __v1__write_req_not_has_been_sent;
  assign __v0__read_req_valid_and_not_has_been_sent = __v0__read_req_vld_buf & __v0__read_req_not_has_been_sent;
  assign __v1__read_req_valid_and_not_has_been_sent = __v0__read_req_vld_buf & __v1__read_req_not_has_been_sent;
  assign __v0__write_req_valid_and_not_has_been_sent = __v0__write_req_vld_buf & __v0__write_req_not_has_been_sent;
  assign y_rd_en__1 = __y__read_req_vld_buf & __y__read_req_not_has_been_sent;
  assign __y__write_req_vld_buf = or_6245 & p1_valid & or_5838;
  assign __y__write_req_not_has_been_sent = ~__y__write_req_has_been_sent_reg;
  assign __out_valid_and_not_has_been_sent = __out_vld_buf & __out_not_has_been_sent;
  assign y_ram_zero_latency0_to_is_not_rdy = ~and_6109;
  assign tuple_index_5845 = y__read_resp_select[31:0];
  assign v0_read_addr = {add_5588, v1_read_addr};
  assign v0_write_addr = and_5516[3:0];
  assign v0_in_select = __for_1_loop_contents_condition ? v0_in : 32'h0000_0000;
  assign v1_write_addr = and_5510[1:0];
  assign v1_in_select = __for_2_loop_contents_condition ? v1_in : 32'h0000_0000;
  assign ____fsm_mv_impl_state__at_most_one_next_value = nor_5593 == one_hot_5607[1] & __fsm_mv_impl_returns_this_activation_vars == one_hot_5607[0];
  assign ____fsm___for_3_loop_state__at_most_one_next_value = nor_5558 == one_hot_5608[1] & __for_4_do_break_with_fsm == one_hot_5608[0];
  assign ____fsm___for_4_loop_state_0__at_most_one_next_value = and_5554 == one_hot_5609[1] & __fsm___for_4_loop_returns_this_activation_vars == one_hot_5609[0];
  assign __fsm_mv_impl_state_2_index = 3'h2;
  assign __fsm_mv_impl_state_3_index = 3'h3;
  assign __fsm_mv_impl_state_4_index = 3'h4;
  assign concat_5565 = {and_5554, __for_5_loop_contents_condition};
  assign y_read_addr__1 = and_5515[1:0];
  assign or_5572 = nor_5558 | __fsm___for_4_loop_returns_this_activation_vars;
  assign concat_6036 = {and_6033, and_6034};
  assign __fsm_mv_impl_state_plus_one = ____fsm_mv_impl_state + __fsm_mv_impl_state_1_index;
  assign v0__read_resp_select = p0_and_5554 ? v0__read_resp : literal_5756;
  assign v1__read_resp_select = p0_and_5554 ? v1__read_resp : literal_5760;
  assign continuation_1_ctx_3__full_condi_output = ~(__this[0] | __this[1]);
  assign __for_1_initial_loop_cond = ~and_5516[4];
  assign __for_2_guarded_update_state_elements = ~(~__fsm_mv_impl_in_state_1 | ~ctx_5__full_condition_continuati_output | and_5510[2]);
  assign __for_3_initial_loop_cond = ~and_5511[5];
  assign __for_4_initial_loop_cond = ~and_5505[5];
  assign __for_5_guarded_update_state_elements = ~(~__fsm_mv_impl_in_state_6 | ~ctx_6__full_condition_continuati_output | and_5515[2]);
  assign concat_6085 = {and_6082, and_6083};
  assign concat_6092 = {and_6089, and_6090};
  assign __v1__write_req_valid_and_all_active_outputs_ready = __v1__write_req_vld_buf & p0_all_active_outputs_ready;
  assign __v1__write_req_valid_and_ready_txfr = __v1__write_req_valid_and_not_has_been_sent & v1__write_req_rdy;
  assign __v0__read_req_valid_and_all_active_outputs_ready = __v0__read_req_vld_buf & p0_all_active_outputs_ready;
  assign __v0__read_req_valid_and_ready_txfr = __v0__read_req_valid_and_not_has_been_sent & v0__read_req_rdy;
  assign __v1__read_req_valid_and_ready_txfr = __v1__read_req_valid_and_not_has_been_sent & v1__read_req_rdy;
  assign __v0__write_req_valid_and_all_active_outputs_ready = __v0__write_req_vld_buf & p0_all_active_outputs_ready;
  assign __v0__write_req_valid_and_ready_txfr = __v0__write_req_valid_and_not_has_been_sent & v0__write_req_rdy;
  assign __y__read_req_valid_and_all_active_outputs_ready = __y__read_req_vld_buf & or_6251;
  assign __y__read_req_valid_and_ready_txfr = y_rd_en__1 & y_ram_zero_latency0_from_skid_rdy;
  assign __y__write_req_valid_and_all_active_outputs_ready = __y__write_req_vld_buf & p2_all_active_outputs_ready;
  assign y_wr_en__1 = __y__write_req_vld_buf & __y__write_req_not_has_been_sent;
  assign __out_valid_and_all_active_outputs_ready = __out_vld_buf & p2_all_active_outputs_ready;
  assign __out_valid_and_ready_txfr = __out_valid_and_not_has_been_sent & out_rdy;
  assign y_ram_zero_latency0_skid_data_load_en = __y_rd_en__1_delay_reg & y_ram_zero_latency0_from_skid_rdy & y_ram_zero_latency0_to_is_not_rdy;
  assign y_ram_zero_latency0_skid_valid_set_zero = __y_ram_zero_latency0_valid_skid_reg & and_6109;
  assign tuple_5733 = {p0_tuple_5586_index0};
  assign tuple_5837 = {{and_5816 | and_5817 | p1_and_5582, and_5816 | and_5818 | p1_and_5583}, y_write_value__5 & {32{p1___fsm___for_4_loop_returns_this_activation_vars}}};
  assign y_read_response__1 = tuple_index_5845 & {32{p1___for_5_loop_contents_condition}};
  assign and_6103 = p1_data_enable & p0_and_5554;
  assign and_6105 = p0_data_enable & __for_1_loop_contents_condition;
  assign and_6108 = p0_data_enable & __for_2_loop_contents_condition;
  assign or_6240 = ~p0_stage_done | ____fsm_mv_impl_state__at_most_one_next_value | rst;
  assign or_6242 = ~p0_stage_done | ____fsm___for_3_loop_state__at_most_one_next_value | rst;
  assign or_6244 = ~p0_stage_done | ____fsm___for_4_loop_state_0__at_most_one_next_value | rst;
  assign p3_enable = 1'h1;
  assign p2_enable = 1'h1;
  assign nand_5851 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & p1___fsm_mv_impl_in_state_1);
  assign nand_5852 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & p1___fsm_mv_impl_in_state_2);
  assign nand_5853 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & p1___fsm_mv_impl_in_state_3);
  assign nand_5854 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & p1___fsm_mv_impl_in_state_4);
  assign smul_5746 = smul32b_32b_x_32b(____fsm___for_4_loop_state_1, ____fsm___for_4_loop_state_2);
  assign __fsm_mv_impl_in_state_2 = ____fsm_mv_impl_state == __fsm_mv_impl_state_2_index;
  assign __fsm_mv_impl_in_state_3 = ____fsm_mv_impl_state == __fsm_mv_impl_state_3_index;
  assign __fsm_mv_impl_in_state_4 = ____fsm_mv_impl_state == __fsm_mv_impl_state_4_index;
  assign not_5663 = ~__fsm___for_4_loop_returns_this_activation_vars;
  assign one_hot_sel_5580 = y_read_addr__1 & {2{concat_5565[0]}} | y_read_addr & {2{concat_5565[1]}};
  assign nand_5664 = ~(__fsm_mv_impl_in_state_6 & ctx_6__full_condition_continuati_output);
  assign nand_5665 = ~(__fsm_mv_impl_in_state_5 & ctx_5__full_condition_ctx_6__ful_output & ~____fsm___for_3_loop_state);
  assign and_5582 = or_5572 & and_5511[1];
  assign and_5583 = or_5572 & and_5511[0];
  assign one_hot_sel_6037 = __fsm_mv_impl_state_0_index & {3{concat_6036[0]}} | __fsm_mv_impl_state_plus_one & {3{concat_6036[1]}};
  assign or_6038 = and_6033 | and_6034;
  assign v0_read_response = v0__read_resp_select[31:0];
  assign and_6052 = p0___fsm___for_4_loop_in_state_0 & p1_data_enable;
  assign v1_read_response = v1__read_resp_select[31:0];
  assign y_read_response = tuple_index_5845 & {32{p1_and_5554}};
  assign and_6058 = p1___fsm___for_4_loop_in_state_0 & p2_stage_done;
  assign and_6061 = __for_5_loop_contents_condition & p0_data_enable;
  assign unexpand_for_this_next__1_case_1 = literal_5421[__this];
  assign unexpand_for___for_1__i_next__1_case_1 = add_5534[4:0];
  assign and_6261 = __fsm_mv_impl_in_state_0 & continuation_1_ctx_3__full_condi_output & __for_1_initial_loop_cond & p0_data_enable;
  assign unexpand_for___for_2__i_next__1_case_1 = add_5527[2:0];
  assign and_6070 = __for_2_guarded_update_state_elements & p0_data_enable;
  assign unexpand_for___for_3_i_next__1_case_1 = add_5528[5:0];
  assign and_6262 = __for_4_do_break_with_fsm & __for_3_initial_loop_cond & p0_data_enable;
  assign unexpand_for___for_4_j_next__1_case_1 = add_5519[5:0];
  assign and_6263 = __fsm___for_4_loop_returns_this_activation_vars & __for_4_initial_loop_cond & p0_data_enable;
  assign unexpand_for___for_5__i_next__1_case_1 = add_5532[2:0];
  assign and_6079 = __for_5_guarded_update_state_elements & p0_data_enable;
  assign one_hot_sel_6086 = __fsm___for_4_loop_default_next_state & concat_6085[0] | __for_4_enter_condition & concat_6085[1];
  assign or_6087 = and_6082 | and_6083;
  assign one_hot_sel_6093 = __fsm___for_4_loop_default_next_state & concat_6092[0] | __for_4_enter_condition & concat_6092[1];
  assign or_6094 = and_6089 | and_6090;
  assign __v1__write_req_not_stage_load = ~__v1__write_req_valid_and_all_active_outputs_ready;
  assign __v1__write_req_has_been_sent_reg_load_en = __v1__write_req_valid_and_ready_txfr | __v1__write_req_valid_and_all_active_outputs_ready;
  assign __v0__read_req_not_stage_load = ~__v0__read_req_valid_and_all_active_outputs_ready;
  assign __v0__read_req_has_been_sent_reg_load_en = __v0__read_req_valid_and_ready_txfr | __v0__read_req_valid_and_all_active_outputs_ready;
  assign __v1__read_req_has_been_sent_reg_load_en = __v1__read_req_valid_and_ready_txfr | __v0__read_req_valid_and_all_active_outputs_ready;
  assign __v0__write_req_not_stage_load = ~__v0__write_req_valid_and_all_active_outputs_ready;
  assign __v0__write_req_has_been_sent_reg_load_en = __v0__write_req_valid_and_ready_txfr | __v0__write_req_valid_and_all_active_outputs_ready;
  assign __y__read_req_not_stage_load = ~__y__read_req_valid_and_all_active_outputs_ready;
  assign __y__read_req_has_been_sent_reg_load_en = __y__read_req_valid_and_ready_txfr | __y__read_req_valid_and_all_active_outputs_ready;
  assign __y__write_req_not_stage_load = ~__y__write_req_valid_and_all_active_outputs_ready;
  assign __y__write_req_has_been_sent_reg_load_en = y_wr_en__1 | __y__write_req_valid_and_all_active_outputs_ready;
  assign __out_not_stage_load = ~__out_valid_and_all_active_outputs_ready;
  assign __out_has_been_sent_reg_load_en = __out_valid_and_ready_txfr | __out_valid_and_all_active_outputs_ready;
  assign y_ram_zero_latency0_skid_valid_load_en = y_ram_zero_latency0_skid_data_load_en | y_ram_zero_latency0_skid_valid_set_zero;
  always_ff @ (posedge clk) begin
    if (rst) begin
      ____for_4__last_iter_broke <= 1'h1;
      ____for_2__last_iter_broke <= 1'h1;
      ____for_3__last_iter_broke <= 1'h1;
      ____for_5__last_iter_broke <= 1'h1;
      ____for_1__last_iter_broke <= 1'h1;
      ____for_4_j <= 6'h00;
      ____for_2__i <= 3'h0;
      ____for_3_i <= 6'h00;
      ____for_5__i <= 3'h0;
      ____for_1__i <= 5'h00;
      ____fsm_mv_impl_state <= 3'h0;
      __this <= 2'h0;
      ____fsm___for_3_loop_state <= 1'h0;
      ____fsm___for_4_loop_state_0 <= 1'h0;
      p0_____fsm___for_4_loop_state_0__1 <= 1'h0;
      p0___fsm_mv_impl_in_state_1 <= 1'h0;
      p0___for_2_loop_contents_condition <= 1'h0;
      p0_ctx_5__full_condition_ctx_6__ful_output <= 1'h0;
      p0___fsm___for_4_loop_in_state_0 <= 1'h0;
      p0___fsm___for_4_loop_returns_this_activation_vars <= 1'h0;
      p0___for_5_loop_contents_condition <= 1'h0;
      p0___fsm_mv_impl_in_state_2 <= 1'h0;
      p0___fsm_mv_impl_in_state_3 <= 1'h0;
      p0___fsm_mv_impl_in_state_4 <= 1'h0;
      p0_and_5554 <= 1'h0;
      p0___for_1_loop_contents_condition <= 1'h0;
      p0_nor_5558 <= 1'h0;
      p0_not_5663 <= 1'h0;
      p0_tuple_5586_index0 <= 2'h0;
      p0_nand_5664 <= 1'h0;
      p0_nand_5665 <= 1'h0;
      p0_and_5582 <= 1'h0;
      p0_and_5583 <= 1'h0;
      ____fsm___for_4_loop_state_1 <= 32'h0000_0000;
      ____fsm___for_4_loop_state_2 <= 32'h0000_0000;
      p1_____fsm___for_4_loop_state_0__1 <= 1'h0;
      p1___fsm_mv_impl_in_state_1 <= 1'h0;
      p1_ctx_5__full_condition_ctx_6__ful_output <= 1'h0;
      p1_smul_5746 <= 32'h0000_0000;
      p1___fsm___for_4_loop_in_state_0 <= 1'h0;
      p1___fsm___for_4_loop_returns_this_activation_vars <= 1'h0;
      p1___for_5_loop_contents_condition <= 1'h0;
      p1___fsm_mv_impl_in_state_2 <= 1'h0;
      p1___fsm_mv_impl_in_state_3 <= 1'h0;
      p1___fsm_mv_impl_in_state_4 <= 1'h0;
      p1_and_5554 <= 1'h0;
      p1_nor_5558 <= 1'h0;
      p1_not_5663 <= 1'h0;
      p1_not_5767 <= 1'h0;
      p1_or_5748 <= 1'h0;
      p1_nand_5664 <= 1'h0;
      p1_nand_5665 <= 1'h0;
      p1_and_5582 <= 1'h0;
      p1_and_5583 <= 1'h0;
      ____fsm___for_4_loop_state_3 <= 32'h0000_0000;
      p2___fsm___for_4_loop_returns_this_activation_vars <= 1'h0;
      p2_nor_5558 <= 1'h0;
      p2_and_5834 <= 1'h0;
      p2_and_5818 <= 1'h0;
      p2_and_5817 <= 1'h0;
      p2_and_5816 <= 1'h0;
      p2_not_5663 <= 1'h0;
      p2_or_5838 <= 1'h0;
      p2_nand_5665 <= 1'h0;
      p2_nand_5851 <= 1'h0;
      p2_nand_5852 <= 1'h0;
      p2_nand_5853 <= 1'h0;
      p2_nand_5854 <= 1'h0;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      __v1__write_req_has_been_sent_reg <= 1'h0;
      __v0__read_req_has_been_sent_reg <= 1'h0;
      __v1__read_req_has_been_sent_reg <= 1'h0;
      __v0__write_req_has_been_sent_reg <= 1'h0;
      __y__read_req_has_been_sent_reg <= 1'h0;
      __y__write_req_has_been_sent_reg <= 1'h0;
      __out_has_been_sent_reg <= 1'h0;
      __y_rd_en__1_delay_reg <= 1'h0;
      __y_ram_zero_latency0_skid_reg <= 32'h0000_0000;
      __y_ram_zero_latency0_valid_skid_reg <= 1'h0;
    end else begin
      ____for_4__last_iter_broke <= and_6090 ? __for_4_do_break_from_func : ____for_4__last_iter_broke;
      ____for_2__last_iter_broke <= and_6108 ? __for_2_do_break_from_func : ____for_2__last_iter_broke;
      ____for_3__last_iter_broke <= and_6083 ? __for_3_do_break_from_func : ____for_3__last_iter_broke;
      ____for_5__last_iter_broke <= and_6061 ? __for_5_do_break_from_func : ____for_5__last_iter_broke;
      ____for_1__last_iter_broke <= and_6105 ? __for_1_do_break_from_func : ____for_1__last_iter_broke;
      ____for_4_j <= and_6263 ? unexpand_for___for_4_j_next__1_case_1 : ____for_4_j;
      ____for_2__i <= and_6070 ? unexpand_for___for_2__i_next__1_case_1 : ____for_2__i;
      ____for_3_i <= and_6262 ? unexpand_for___for_3_i_next__1_case_1 : ____for_3_i;
      ____for_5__i <= and_6079 ? unexpand_for___for_5__i_next__1_case_1 : ____for_5__i;
      ____for_1__i <= and_6261 ? unexpand_for___for_1__i_next__1_case_1 : ____for_1__i;
      ____fsm_mv_impl_state <= or_6038 ? one_hot_sel_6037 : ____fsm_mv_impl_state;
      __this <= and_6034 ? unexpand_for_this_next__1_case_1 : __this;
      ____fsm___for_3_loop_state <= or_6087 ? one_hot_sel_6086 : ____fsm___for_3_loop_state;
      ____fsm___for_4_loop_state_0 <= or_6094 ? one_hot_sel_6093 : ____fsm___for_4_loop_state_0;
      p0_____fsm___for_4_loop_state_0__1 <= p0_data_enable ? ____fsm___for_4_loop_state_0 : p0_____fsm___for_4_loop_state_0__1;
      p0___fsm_mv_impl_in_state_1 <= p0_data_enable ? __fsm_mv_impl_in_state_1 : p0___fsm_mv_impl_in_state_1;
      p0___for_2_loop_contents_condition <= p0_data_enable ? __for_2_loop_contents_condition : p0___for_2_loop_contents_condition;
      p0_ctx_5__full_condition_ctx_6__ful_output <= p0_data_enable ? ctx_5__full_condition_ctx_6__ful_output : p0_ctx_5__full_condition_ctx_6__ful_output;
      p0___fsm___for_4_loop_in_state_0 <= p0_data_enable ? __fsm___for_4_loop_in_state_0 : p0___fsm___for_4_loop_in_state_0;
      p0___fsm___for_4_loop_returns_this_activation_vars <= p0_data_enable ? __fsm___for_4_loop_returns_this_activation_vars : p0___fsm___for_4_loop_returns_this_activation_vars;
      p0___for_5_loop_contents_condition <= p0_data_enable ? __for_5_loop_contents_condition : p0___for_5_loop_contents_condition;
      p0___fsm_mv_impl_in_state_2 <= p0_data_enable ? __fsm_mv_impl_in_state_2 : p0___fsm_mv_impl_in_state_2;
      p0___fsm_mv_impl_in_state_3 <= p0_data_enable ? __fsm_mv_impl_in_state_3 : p0___fsm_mv_impl_in_state_3;
      p0___fsm_mv_impl_in_state_4 <= p0_data_enable ? __fsm_mv_impl_in_state_4 : p0___fsm_mv_impl_in_state_4;
      p0_and_5554 <= p0_data_enable ? and_5554 : p0_and_5554;
      p0___for_1_loop_contents_condition <= p0_data_enable ? __for_1_loop_contents_condition : p0___for_1_loop_contents_condition;
      p0_nor_5558 <= p0_data_enable ? nor_5558 : p0_nor_5558;
      p0_not_5663 <= p0_data_enable ? not_5663 : p0_not_5663;
      p0_tuple_5586_index0 <= p0_data_enable ? one_hot_sel_5580 : p0_tuple_5586_index0;
      p0_nand_5664 <= p0_data_enable ? nand_5664 : p0_nand_5664;
      p0_nand_5665 <= p0_data_enable ? nand_5665 : p0_nand_5665;
      p0_and_5582 <= p0_data_enable ? and_5582 : p0_and_5582;
      p0_and_5583 <= p0_data_enable ? and_5583 : p0_and_5583;
      ____fsm___for_4_loop_state_1 <= and_6052 ? v0_read_response : ____fsm___for_4_loop_state_1;
      ____fsm___for_4_loop_state_2 <= and_6052 ? v1_read_response : ____fsm___for_4_loop_state_2;
      p1_____fsm___for_4_loop_state_0__1 <= p1_data_enable ? p0_____fsm___for_4_loop_state_0__1 : p1_____fsm___for_4_loop_state_0__1;
      p1___fsm_mv_impl_in_state_1 <= p1_data_enable ? p0___fsm_mv_impl_in_state_1 : p1___fsm_mv_impl_in_state_1;
      p1_ctx_5__full_condition_ctx_6__ful_output <= p1_data_enable ? p0_ctx_5__full_condition_ctx_6__ful_output : p1_ctx_5__full_condition_ctx_6__ful_output;
      p1_smul_5746 <= p1_data_enable ? smul_5746 : p1_smul_5746;
      p1___fsm___for_4_loop_in_state_0 <= p1_data_enable ? p0___fsm___for_4_loop_in_state_0 : p1___fsm___for_4_loop_in_state_0;
      p1___fsm___for_4_loop_returns_this_activation_vars <= p1_data_enable ? p0___fsm___for_4_loop_returns_this_activation_vars : p1___fsm___for_4_loop_returns_this_activation_vars;
      p1___for_5_loop_contents_condition <= p1_data_enable ? p0___for_5_loop_contents_condition : p1___for_5_loop_contents_condition;
      p1___fsm_mv_impl_in_state_2 <= p1_data_enable ? p0___fsm_mv_impl_in_state_2 : p1___fsm_mv_impl_in_state_2;
      p1___fsm_mv_impl_in_state_3 <= p1_data_enable ? p0___fsm_mv_impl_in_state_3 : p1___fsm_mv_impl_in_state_3;
      p1___fsm_mv_impl_in_state_4 <= p1_data_enable ? p0___fsm_mv_impl_in_state_4 : p1___fsm_mv_impl_in_state_4;
      p1_and_5554 <= p1_data_enable ? p0_and_5554 : p1_and_5554;
      p1_nor_5558 <= p1_data_enable ? p0_nor_5558 : p1_nor_5558;
      p1_not_5663 <= p1_data_enable ? p0_not_5663 : p1_not_5663;
      p1_not_5767 <= p1_data_enable ? not_5904 : p1_not_5767;
      p1_or_5748 <= p1_data_enable ? or_5748 : p1_or_5748;
      p1_nand_5664 <= p1_data_enable ? p0_nand_5664 : p1_nand_5664;
      p1_nand_5665 <= p1_data_enable ? p0_nand_5665 : p1_nand_5665;
      p1_and_5582 <= p1_data_enable ? p0_and_5582 : p1_and_5582;
      p1_and_5583 <= p1_data_enable ? p0_and_5583 : p1_and_5583;
      ____fsm___for_4_loop_state_3 <= and_6058 ? y_read_response : ____fsm___for_4_loop_state_3;
      p2___fsm___for_4_loop_returns_this_activation_vars <= p2_stage_done ? p1___fsm___for_4_loop_returns_this_activation_vars : p2___fsm___for_4_loop_returns_this_activation_vars;
      p2_nor_5558 <= p2_stage_done ? p1_nor_5558 : p2_nor_5558;
      p2_and_5834 <= p2_stage_done ? and_5834 : p2_and_5834;
      p2_and_5818 <= p2_stage_done ? and_5818 : p2_and_5818;
      p2_and_5817 <= p2_stage_done ? and_5817 : p2_and_5817;
      p2_and_5816 <= p2_stage_done ? and_5816 : p2_and_5816;
      p2_not_5663 <= p2_stage_done ? p1_not_5663 : p2_not_5663;
      p2_or_5838 <= p2_stage_done ? or_5838 : p2_or_5838;
      p2_nand_5665 <= p2_stage_done ? p1_nand_5665 : p2_nand_5665;
      p2_nand_5851 <= p2_stage_done ? nand_5851 : p2_nand_5851;
      p2_nand_5852 <= p2_stage_done ? nand_5852 : p2_nand_5852;
      p2_nand_5853 <= p2_stage_done ? nand_5853 : p2_nand_5853;
      p2_nand_5854 <= p2_stage_done ? nand_5854 : p2_nand_5854;
      p0_valid <= p0_enable ? p0_stage_done : p0_valid;
      p1_valid <= p1_enable ? p1_stage_done : p1_valid;
      p2_valid <= p2_enable ? p2_stage_done : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      __v1__write_req_has_been_sent_reg <= __v1__write_req_has_been_sent_reg_load_en ? __v1__write_req_not_stage_load : __v1__write_req_has_been_sent_reg;
      __v0__read_req_has_been_sent_reg <= __v0__read_req_has_been_sent_reg_load_en ? __v0__read_req_not_stage_load : __v0__read_req_has_been_sent_reg;
      __v1__read_req_has_been_sent_reg <= __v1__read_req_has_been_sent_reg_load_en ? __v0__read_req_not_stage_load : __v1__read_req_has_been_sent_reg;
      __v0__write_req_has_been_sent_reg <= __v0__write_req_has_been_sent_reg_load_en ? __v0__write_req_not_stage_load : __v0__write_req_has_been_sent_reg;
      __y__read_req_has_been_sent_reg <= __y__read_req_has_been_sent_reg_load_en ? __y__read_req_not_stage_load : __y__read_req_has_been_sent_reg;
      __y__write_req_has_been_sent_reg <= __y__write_req_has_been_sent_reg_load_en ? __y__write_req_not_stage_load : __y__write_req_has_been_sent_reg;
      __out_has_been_sent_reg <= __out_has_been_sent_reg_load_en ? __out_not_stage_load : __out_has_been_sent_reg;
      __y_rd_en__1_delay_reg <= y_rd_en__1;
      __y_ram_zero_latency0_skid_reg <= y_ram_zero_latency0_skid_data_load_en ? y_rd_data : __y_ram_zero_latency0_skid_reg;
      __y_ram_zero_latency0_valid_skid_reg <= y_ram_zero_latency0_skid_valid_load_en ? y_ram_zero_latency0_from_skid_rdy : __y_ram_zero_latency0_valid_skid_reg;
    end
  end
  assign out = y_read_response__1;
  assign out_vld = __out_valid_and_not_has_been_sent;
  assign v0__read_req = {v0_read_addr};
  assign v0__read_req_vld = __v0__read_req_valid_and_not_has_been_sent;
  assign v0__read_resp_rdy = and_6103;
  assign v0__write_completion_rdy = p1_data_enable & p0___for_1_loop_contents_condition;
  assign v0__write_req = {v0_write_addr, v0_in_select};
  assign v0__write_req_vld = __v0__write_req_valid_and_not_has_been_sent;
  assign v0_in_rdy = and_6105;
  assign v1__read_req = {v1_read_addr};
  assign v1__read_req_vld = __v1__read_req_valid_and_not_has_been_sent;
  assign v1__read_resp_rdy = and_6103;
  assign v1__write_completion_rdy = p1_data_enable & p0___for_2_loop_contents_condition;
  assign v1__write_req = {v1_write_addr, v1_in_select};
  assign v1__write_req_vld = __v1__write_req_valid_and_not_has_been_sent;
  assign v1_in_rdy = and_6108;
  assign y_rd_addr = tuple_5733[1:0];
  assign y_rd_en = y_rd_en__1;
  assign y_wr_addr = tuple_5837[33:32];
  assign y_wr_data = tuple_5837[31:0];
  assign y_wr_en = y_wr_en__1;
  `ifdef ASSERT_ON
  ____fsm_mv_impl_state__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_6240))) or_6240) else $fatal(0, "More than one next_value fired for state element: __fsm_mv_impl_state");
  ____fsm___for_3_loop_state__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_6242))) or_6242) else $fatal(0, "More than one next_value fired for state element: __fsm___for_3_loop_state");
  ____fsm___for_4_loop_state_0__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_6244))) or_6244) else $fatal(0, "More than one next_value fired for state element: __fsm___for_4_loop_state_0");
  `endif  // ASSERT_ON
endmodule