module gemm_mem(
  input wire clk,
  input wire rst,
  input wire out_rdy,
  input wire v0__read_req_rdy,
  input wire [31:0] v0__read_resp,
  input wire v0__read_resp_vld,
  input wire v0__write_completion_vld,
  input wire v0__write_req_rdy,
  input wire [31:0] v0_in,
  input wire v0_in_vld,
  input wire v1__read_req_rdy,
  input wire [31:0] v1__read_resp,
  input wire v1__read_resp_vld,
  input wire v1__write_completion_vld,
  input wire v1__write_req_rdy,
  input wire [31:0] v1_in,
  input wire v1_in_vld,
  input wire [31:0] C_rd_data,
  output wire [31:0] out,
  output wire out_vld,
  output wire [3:0] v0__read_req,
  output wire v0__read_req_vld,
  output wire v0__read_resp_rdy,
  output wire v0__write_completion_rdy,
  output wire [35:0] v0__write_req,
  output wire v0__write_req_vld,
  output wire v0_in_rdy,
  output wire [3:0] v1__read_req,
  output wire v1__read_req_vld,
  output wire v1__read_resp_rdy,
  output wire v1__write_completion_rdy,
  output wire [35:0] v1__write_req,
  output wire v1__write_req_vld,
  output wire v1_in_rdy,
  output wire [3:0] C_rd_addr,
  output wire C_rd_en,
  output wire [3:0] C_wr_addr,
  output wire [31:0] C_wr_data,
  output wire C_wr_en
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] smul32b_32b_x_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    reg signed [31:0] signed_lhs;
    reg signed [31:0] signed_rhs;
    reg signed [31:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul32b_32b_x_32b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  wire [31:0] literal_11959 = 32'h0000_0000;
  wire [31:0] literal_11836 = 32'h0000_0000;
  wire [31:0] literal_11840 = 32'h0000_0000;
  wire [1:0] literal_11493[4];
  assign literal_11493 = '{2'h1, 2'h2, 2'h3, 2'h0};
  reg ____for_5__last_iter_broke;
  reg ____for_4__last_iter_broke;
  reg ____for_2__last_iter_broke;
  reg ____for_3__last_iter_broke;
  reg [2:0] ____for_5_k;
  reg ____for_6__last_iter_broke;
  reg ____for_1__last_iter_broke;
  reg [2:0] ____for_4_j;
  reg [4:0] ____for_2__i;
  reg [2:0] ____for_3_i;
  reg [1:0] __this;
  reg [4:0] ____for_6__i;
  reg [4:0] ____for_1__i;
  reg [4:0] ____fsm_gemm_impl_state;
  reg ____fsm___for_5_loop_state_0;
  reg [4:0] p0_____fsm_gemm_impl_state__1;
  reg p0_____fsm___for_5_loop_state_0__1;
  reg p0___fsm_gemm_impl_in_state_1;
  reg p0___for_2_loop_contents_condition;
  reg p0_ctx_5__full_condition_ctx_6__ful_output;
  reg p0___fsm___for_5_loop_in_state_0;
  reg p0___fsm___for_5_loop_returns_this_activation_vars;
  reg p0___for_6_loop_contents_condition;
  reg p0_nor_11636;
  reg p0___for_1_loop_contents_condition;
  reg [3:0] p0_tuple_11671_index0;
  reg p0_nand_11745;
  reg p0_nand_11746;
  reg p0_nand_11747;
  reg p0_and_11664;
  reg p0_and_11665;
  reg p0_and_11666;
  reg p0_and_11667;
  reg [31:0] ____fsm___for_5_loop_state_1;
  reg [31:0] ____fsm___for_5_loop_state_2;
  reg [4:0] p1_____fsm_gemm_impl_state__1;
  reg p1_____fsm___for_5_loop_state_0__1;
  reg p1___fsm_gemm_impl_in_state_1;
  reg p1_ctx_5__full_condition_ctx_6__ful_output;
  reg p1___fsm___for_5_loop_in_state_0;
  reg p1___fsm___for_5_loop_returns_this_activation_vars;
  reg [31:0] p1_smul_11826;
  reg p1___for_6_loop_contents_condition;
  reg p1_nor_11636;
  reg p1_or_11828;
  reg p1_nand_11745;
  reg p1_nand_11746;
  reg p1_nand_11747;
  reg p1_and_11664;
  reg p1_and_11665;
  reg p1_and_11666;
  reg p1_and_11667;
  reg [31:0] ____fsm___for_5_loop_state_3;
  reg p2___fsm___for_5_loop_returns_this_activation_vars;
  reg p2_and_11953;
  reg p2_and_11924;
  reg p2_and_11923;
  reg p2_and_11912;
  reg p2_and_11921;
  reg p2_and_11908;
  reg p2_and_11906;
  reg p2_and_11898;
  reg p2_and_11918;
  reg p2_and_11917;
  reg p2_and_11916;
  reg p2_and_11911;
  reg p2_and_11915;
  reg p2_and_11907;
  reg p2_and_11905;
  reg p2_and_11897;
  reg p2_or_11957;
  reg p2_nand_11745;
  reg p2_nand_11970;
  reg p2_nand_11971;
  reg p2_nand_11972;
  reg p2_nand_11973;
  reg p2_nand_11974;
  reg p2_nand_11975;
  reg p2_nand_11976;
  reg p2_nand_11977;
  reg p2_nand_11978;
  reg p2_nand_11979;
  reg p2_nand_11980;
  reg p2_nand_11981;
  reg p2_nand_11982;
  reg p2_nand_11983;
  reg p2_nand_11984;
  reg p2_nand_11985;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg __v1__write_req_has_been_sent_reg;
  reg __v0__read_req_has_been_sent_reg;
  reg __v1__read_req_has_been_sent_reg;
  reg __v0__write_req_has_been_sent_reg;
  reg __C__read_req_has_been_sent_reg;
  reg __C__write_req_has_been_sent_reg;
  reg __out_has_been_sent_reg;
  reg __C_rd_en__1_delay_reg;
  reg [31:0] __C_ram_zero_latency0_skid_reg;
  reg __C_ram_zero_latency0_valid_skid_reg;
  wire __fsm___for_5_loop_default_next_state;
  wire [2:0] and_11575;
  wire [2:0] and_11582;
  wire [4:0] and_11589;
  wire [2:0] and_11590;
  wire [3:0] add_11592;
  wire [4:0] __fsm_gemm_impl_state_17_index;
  wire ctx_5__full_condition_ctx_6__ful_output;
  wire [4:0] and_11596;
  wire [4:0] and_11597;
  wire [3:0] add_11600;
  wire [1:0] __fsm___for_5_loop_initial_state_index;
  wire ne_11602;
  wire __for_3_not_enter_condition;
  wire __fsm___for_5_loop_in_state_0;
  wire [5:0] add_11609;
  wire [3:0] add_11610;
  wire __for_5_do_break_from_func;
  wire __fsm___for_5_loop_returns_this_activation_vars;
  wire [5:0] add_11614;
  wire [5:0] add_11617;
  wire __for_4_do_break_from_func;
  wire __for_5_do_break_with_fsm;
  wire __for_2_do_break_from_func;
  wire __for_3_do_break_from_func;
  wire __for_4_do_break_with_fsm;
  wire __for_6_do_break_from_func;
  wire [4:0] __fsm_gemm_impl_state_0_index;
  wire __for_1_do_break_from_func;
  wire ctx_5__full_condition_continuati_output;
  wire __for_3_do_break_with_fsm;
  wire ctx_6__full_condition_continuati_output;
  wire [4:0] __fsm_gemm_impl_state_1_index;
  wire __fsm_gemm_impl_in_state_0;
  wire __for_1_not_exit_state_condition;
  wire __for_2_not_exit_state_condition;
  wire __for_4_enter_condition;
  wire __for_3_not_exit_state_condition;
  wire __for_6_not_exit_state_condition;
  wire or_11828;
  wire __fsm_gemm_impl_in_state_1;
  wire __fsm_gemm_impl_go_to_next_state_in_state;
  wire [4:0] __fsm_gemm_impl_state_18_index;
  wire or_12447;
  wire p2_all_active_outputs_ready;
  wire C__read_req_not_pred;
  wire C_ram_zero_latency0_from_skid_rdy;
  wire __for_2_loop_contents_condition;
  wire __for_1_loop_contents_condition;
  wire nor_11636;
  wire [4:0] __fsm_gemm_impl_state_16_index;
  wire [4:0] __fsm_gemm_impl_state_8_index;
  wire __fsm_gemm_impl_in_state_18;
  wire p2_stage_done;
  wire p2_not_valid;
  wire p1_all_active_inputs_valid;
  wire or_12453;
  wire v0__read_req_not_pred;
  wire [4:0] __fsm_gemm_impl_state_15_index;
  wire [4:0] __fsm_gemm_impl_state_7_index;
  wire [4:0] __fsm_gemm_impl_state_14_index;
  wire [4:0] __fsm_gemm_impl_state_6_index;
  wire __fsm_gemm_impl_in_state_16;
  wire __fsm_gemm_impl_in_state_8;
  wire [4:0] __fsm_gemm_impl_state_12_index;
  wire [4:0] __fsm_gemm_impl_state_4_index;
  wire nor_11679;
  wire __fsm_gemm_impl_returns_this_activation_vars;
  wire p1_enable;
  wire p1_stage_done;
  wire [4:0] __fsm_gemm_impl_state_2_index;
  wire [4:0] __fsm_gemm_impl_state_3_index;
  wire [4:0] __fsm_gemm_impl_state_5_index;
  wire [4:0] __fsm_gemm_impl_state_9_index;
  wire [4:0] __fsm_gemm_impl_state_10_index;
  wire [4:0] __fsm_gemm_impl_state_11_index;
  wire [4:0] __fsm_gemm_impl_state_13_index;
  wire __fsm_gemm_impl_in_state_15;
  wire __fsm_gemm_impl_in_state_7;
  wire __fsm_gemm_impl_in_state_14;
  wire __fsm_gemm_impl_in_state_6;
  wire and_11897;
  wire and_11898;
  wire __fsm_gemm_impl_in_state_12;
  wire __fsm_gemm_impl_in_state_4;
  wire [1:0] ____fsm_gemm_impl_state__next_value_predicates;
  wire [1:0] ____fsm___for_5_loop_state_0__next_value_predicates;
  wire p1_data_enable;
  wire p1_not_valid;
  wire p0_all_active_inputs_valid;
  wire p0_all_active_outputs_ready;
  wire __fsm_gemm_impl_in_state_2;
  wire __fsm_gemm_impl_in_state_3;
  wire __fsm_gemm_impl_in_state_5;
  wire __fsm_gemm_impl_in_state_9;
  wire __fsm_gemm_impl_in_state_10;
  wire __fsm_gemm_impl_in_state_11;
  wire __fsm_gemm_impl_in_state_13;
  wire and_11905;
  wire and_11906;
  wire and_11907;
  wire and_11908;
  wire or_11910;
  wire and_11911;
  wire and_11912;
  wire [31:0] C_ram_zero_latency0_select;
  wire [2:0] one_hot_11692;
  wire [2:0] one_hot_11693;
  wire p0_enable;
  wire p0_stage_done;
  wire and_11953;
  wire and_11924;
  wire and_11923;
  wire and_11921;
  wire and_11918;
  wire and_11917;
  wire and_11916;
  wire and_11915;
  wire or_11919;
  wire or_11920;
  wire or_11922;
  wire [1:0] concat_11626;
  wire p0_data_enable;
  wire __v1__write_req_vld_buf;
  wire __v1__write_req_not_has_been_sent;
  wire __v0__read_req_vld_buf;
  wire __v0__read_req_not_has_been_sent;
  wire __v1__read_req_not_has_been_sent;
  wire __v0__write_req_vld_buf;
  wire __v0__write_req_not_has_been_sent;
  wire __C__read_req_vld_buf;
  wire __C__read_req_not_has_been_sent;
  wire or_11957;
  wire __out_vld_buf;
  wire __out_not_has_been_sent;
  wire and_12307;
  wire [31:0] C_write_value__16;
  wire [31:0] C__read_resp_select;
  wire [1:0] add_11673;
  wire [1:0] add_11674;
  wire __for_6_loop_contents_condition;
  wire [1:0] add_11638;
  wire and_12238;
  wire and_12239;
  wire and_12293;
  wire and_12294;
  wire __v1__write_req_valid_and_not_has_been_sent;
  wire __v0__read_req_valid_and_not_has_been_sent;
  wire __v1__read_req_valid_and_not_has_been_sent;
  wire __v0__write_req_valid_and_not_has_been_sent;
  wire C_rd_en__1;
  wire __C__write_req_vld_buf;
  wire __C__write_req_not_has_been_sent;
  wire __out_valid_and_not_has_been_sent;
  wire C_ram_zero_latency0_to_is_not_rdy;
  wire [31:0] tuple_index_11964;
  wire [3:0] v0_read_addr;
  wire [3:0] v0_write_addr;
  wire [31:0] v0_in_select;
  wire [3:0] v1_read_addr;
  wire [3:0] v1_write_addr;
  wire [31:0] v1_in_select;
  wire ____fsm_gemm_impl_state__at_most_one_next_value;
  wire ____fsm___for_5_loop_state_0__at_most_one_next_value;
  wire [1:0] concat_11648;
  wire [3:0] C_read_addr__1;
  wire [3:0] C_read_addr;
  wire [1:0] concat_12241;
  wire [4:0] __fsm_gemm_impl_state_plus_one;
  wire [31:0] v0__read_resp_select;
  wire [31:0] v1__read_resp_select;
  wire continuation_1_ctx_3__full_condi_output;
  wire __for_1_initial_loop_cond;
  wire __for_2_guarded_update_state_elements;
  wire __for_3_initial_loop_cond;
  wire __for_4_initial_loop_cond;
  wire __for_5_initial_loop_cond;
  wire __for_6_guarded_update_state_elements;
  wire [1:0] concat_12296;
  wire __v1__write_req_valid_and_all_active_outputs_ready;
  wire __v1__write_req_valid_and_ready_txfr;
  wire __v0__read_req_valid_and_all_active_outputs_ready;
  wire __v0__read_req_valid_and_ready_txfr;
  wire __v1__read_req_valid_and_ready_txfr;
  wire __v0__write_req_valid_and_all_active_outputs_ready;
  wire __v0__write_req_valid_and_ready_txfr;
  wire __C__read_req_valid_and_all_active_outputs_ready;
  wire __C__read_req_valid_and_ready_txfr;
  wire __C__write_req_valid_and_all_active_outputs_ready;
  wire C_wr_en__1;
  wire __out_valid_and_all_active_outputs_ready;
  wire __out_valid_and_ready_txfr;
  wire C_ram_zero_latency0_skid_data_load_en;
  wire C_ram_zero_latency0_skid_valid_set_zero;
  wire [3:0] tuple_11807;
  wire [35:0] tuple_11956;
  wire [31:0] C_read_response__1;
  wire and_12309;
  wire and_12311;
  wire and_12314;
  wire or_12444;
  wire or_12446;
  wire p3_enable;
  wire p2_enable;
  wire nand_11970;
  wire nand_11971;
  wire nand_11972;
  wire nand_11973;
  wire nand_11974;
  wire nand_11975;
  wire nand_11976;
  wire nand_11977;
  wire nand_11978;
  wire nand_11979;
  wire nand_11980;
  wire nand_11981;
  wire nand_11982;
  wire nand_11983;
  wire nand_11984;
  wire nand_11985;
  wire [31:0] smul_11826;
  wire [3:0] one_hot_sel_11662;
  wire nand_11745;
  wire nand_11746;
  wire nand_11747;
  wire and_11664;
  wire and_11665;
  wire and_11666;
  wire and_11667;
  wire [4:0] one_hot_sel_12242;
  wire or_12243;
  wire and_12251;
  wire and_12254;
  wire [31:0] v0_read_response;
  wire and_12260;
  wire [31:0] v1_read_response;
  wire [31:0] C_read_response;
  wire and_12266;
  wire and_12269;
  wire [1:0] unexpand_for_this_next__1_case_1;
  wire [4:0] unexpand_for___for_1__i_next__1_case_1;
  wire and_12463;
  wire [4:0] unexpand_for___for_2__i_next__1_case_1;
  wire and_12278;
  wire [2:0] unexpand_for___for_3_i_next__1_case_1;
  wire and_12464;
  wire [2:0] unexpand_for___for_4_j_next__1_case_1;
  wire and_12465;
  wire [2:0] unexpand_for___for_5_k_next__1_case_1;
  wire and_12466;
  wire [4:0] unexpand_for___for_6__i_next__1_case_1;
  wire and_12290;
  wire one_hot_sel_12297;
  wire or_12298;
  wire __v1__write_req_not_stage_load;
  wire __v1__write_req_has_been_sent_reg_load_en;
  wire __v0__read_req_not_stage_load;
  wire __v0__read_req_has_been_sent_reg_load_en;
  wire __v1__read_req_has_been_sent_reg_load_en;
  wire __v0__write_req_not_stage_load;
  wire __v0__write_req_has_been_sent_reg_load_en;
  wire __C__read_req_not_stage_load;
  wire __C__read_req_has_been_sent_reg_load_en;
  wire __C__write_req_not_stage_load;
  wire __C__write_req_has_been_sent_reg_load_en;
  wire __out_not_stage_load;
  wire __out_has_been_sent_reg_load_en;
  wire C_ram_zero_latency0_skid_valid_load_en;
  assign __fsm___for_5_loop_default_next_state = 1'h0;
  assign and_11575 = {3{~____for_5__last_iter_broke}} & ____for_5_k;
  assign and_11582 = {3{~____for_4__last_iter_broke}} & ____for_4_j;
  assign and_11589 = {5{~____for_2__last_iter_broke}} & ____for_2__i;
  assign and_11590 = {3{~____for_3__last_iter_broke}} & ____for_3_i;
  assign add_11592 = {__fsm___for_5_loop_default_next_state, and_11575} + 4'h1;
  assign __fsm_gemm_impl_state_17_index = 5'h11;
  assign ctx_5__full_condition_ctx_6__ful_output = __this == 2'h2;
  assign and_11596 = {5{~____for_6__last_iter_broke}} & ____for_6__i;
  assign and_11597 = {5{~____for_1__last_iter_broke}} & ____for_1__i;
  assign add_11600 = {__fsm___for_5_loop_default_next_state, and_11582} + 4'h1;
  assign __fsm___for_5_loop_initial_state_index = 2'h0;
  assign ne_11602 = ____fsm_gemm_impl_state != __fsm_gemm_impl_state_17_index;
  assign __for_3_not_enter_condition = ~ctx_5__full_condition_ctx_6__ful_output;
  assign __fsm___for_5_loop_in_state_0 = ~____fsm___for_5_loop_state_0;
  assign add_11609 = {__fsm___for_5_loop_default_next_state, and_11589} + 6'h01;
  assign add_11610 = {__fsm___for_5_loop_default_next_state, and_11590} + 4'h1;
  assign __for_5_do_break_from_func = add_11592[3:2] != __fsm___for_5_loop_initial_state_index;
  assign __fsm___for_5_loop_returns_this_activation_vars = ~(ne_11602 | __for_3_not_enter_condition | __fsm___for_5_loop_in_state_0);
  assign add_11614 = {__fsm___for_5_loop_default_next_state, and_11596} + 6'h01;
  assign add_11617 = {__fsm___for_5_loop_default_next_state, and_11597} + 6'h01;
  assign __for_4_do_break_from_func = add_11600[3:2] != __fsm___for_5_loop_initial_state_index;
  assign __for_5_do_break_with_fsm = __for_5_do_break_from_func & __fsm___for_5_loop_returns_this_activation_vars;
  assign __for_2_do_break_from_func = add_11609[5:4] != __fsm___for_5_loop_initial_state_index;
  assign __for_3_do_break_from_func = add_11610[3:2] != __fsm___for_5_loop_initial_state_index;
  assign __for_4_do_break_with_fsm = __for_4_do_break_from_func & __for_5_do_break_with_fsm;
  assign __for_6_do_break_from_func = add_11614[5:4] != __fsm___for_5_loop_initial_state_index;
  assign __fsm_gemm_impl_state_0_index = 5'h00;
  assign __for_1_do_break_from_func = add_11617[5:4] != __fsm___for_5_loop_initial_state_index;
  assign ctx_5__full_condition_continuati_output = __this == 2'h1;
  assign __for_3_do_break_with_fsm = __for_3_do_break_from_func & __for_4_do_break_with_fsm;
  assign ctx_6__full_condition_continuati_output = __this == 2'h3;
  assign __fsm_gemm_impl_state_1_index = 5'h01;
  assign __fsm_gemm_impl_in_state_0 = ____fsm_gemm_impl_state == __fsm_gemm_impl_state_0_index;
  assign __for_1_not_exit_state_condition = __this[0] | __this[1] | __for_1_do_break_from_func;
  assign __for_2_not_exit_state_condition = ~(ctx_5__full_condition_continuati_output & ~__for_2_do_break_from_func);
  assign __for_4_enter_condition = 1'h1;
  assign __for_3_not_exit_state_condition = __for_3_not_enter_condition | __for_3_do_break_with_fsm;
  assign __for_6_not_exit_state_condition = ~(ctx_6__full_condition_continuati_output & ~__for_6_do_break_from_func);
  assign or_11828 = p0_nor_11636 | p0___for_6_loop_contents_condition;
  assign __fsm_gemm_impl_in_state_1 = ____fsm_gemm_impl_state == __fsm_gemm_impl_state_1_index;
  assign __fsm_gemm_impl_go_to_next_state_in_state = ____fsm_gemm_impl_state == 5'h00 ? __for_1_not_exit_state_condition : (____fsm_gemm_impl_state == 5'h01 ? __for_2_not_exit_state_condition : (____fsm_gemm_impl_state == 5'h02 ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h03 ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h04 ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h05 ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h06 ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h07 ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h08 ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h09 ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h0a ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h0b ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h0c ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h0d ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h0e ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h0f ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h10 ? __for_4_enter_condition : (____fsm_gemm_impl_state == 5'h11 ? __for_3_not_exit_state_condition : (____fsm_gemm_impl_state == 5'h12 ? __for_6_not_exit_state_condition : __fsm___for_5_loop_default_next_state))))))))))))))))));
  assign __fsm_gemm_impl_state_18_index = 5'h12;
  assign or_12447 = ~p1_or_11828 | __C_rd_en__1_delay_reg | __C_ram_zero_latency0_valid_skid_reg;
  assign p2_all_active_outputs_ready = ~p1___for_6_loop_contents_condition | out_rdy | __out_has_been_sent_reg;
  assign C__read_req_not_pred = ~or_11828;
  assign C_ram_zero_latency0_from_skid_rdy = ~__C_ram_zero_latency0_valid_skid_reg;
  assign __for_2_loop_contents_condition = __fsm_gemm_impl_in_state_1 & ctx_5__full_condition_continuati_output;
  assign __for_1_loop_contents_condition = ~(~__fsm_gemm_impl_in_state_0 | __this[0] | __this[1]);
  assign nor_11636 = ~(ne_11602 | __for_3_not_enter_condition | ____fsm___for_5_loop_state_0);
  assign __fsm_gemm_impl_state_16_index = 5'h10;
  assign __fsm_gemm_impl_state_8_index = 5'h08;
  assign __fsm_gemm_impl_in_state_18 = ____fsm_gemm_impl_state == __fsm_gemm_impl_state_18_index;
  assign p2_stage_done = p1_valid & or_12447 & p2_all_active_outputs_ready;
  assign p2_not_valid = ~p1_valid;
  assign p1_all_active_inputs_valid = (~p0___for_2_loop_contents_condition | v1__write_completion_vld) & (~p0_nor_11636 | v0__read_resp_vld) & (~p0_nor_11636 | v1__read_resp_vld) & (~p0___for_1_loop_contents_condition | v0__write_completion_vld);
  assign or_12453 = C__read_req_not_pred | C_ram_zero_latency0_from_skid_rdy | __C__read_req_has_been_sent_reg;
  assign v0__read_req_not_pred = ~nor_11636;
  assign __fsm_gemm_impl_state_15_index = 5'h0f;
  assign __fsm_gemm_impl_state_7_index = 5'h07;
  assign __fsm_gemm_impl_state_14_index = 5'h0e;
  assign __fsm_gemm_impl_state_6_index = 5'h06;
  assign __fsm_gemm_impl_in_state_16 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_16_index;
  assign __fsm_gemm_impl_in_state_8 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_8_index;
  assign __fsm_gemm_impl_state_12_index = 5'h0c;
  assign __fsm_gemm_impl_state_4_index = 5'h04;
  assign nor_11679 = ~(~__fsm_gemm_impl_go_to_next_state_in_state | __fsm_gemm_impl_in_state_18);
  assign __fsm_gemm_impl_returns_this_activation_vars = __fsm_gemm_impl_in_state_18 & __fsm_gemm_impl_go_to_next_state_in_state;
  assign p1_enable = p2_stage_done | p2_not_valid;
  assign p1_stage_done = p0_valid & p1_all_active_inputs_valid & or_12453;
  assign __fsm_gemm_impl_state_2_index = 5'h02;
  assign __fsm_gemm_impl_state_3_index = 5'h03;
  assign __fsm_gemm_impl_state_5_index = 5'h05;
  assign __fsm_gemm_impl_state_9_index = 5'h09;
  assign __fsm_gemm_impl_state_10_index = 5'h0a;
  assign __fsm_gemm_impl_state_11_index = 5'h0b;
  assign __fsm_gemm_impl_state_13_index = 5'h0d;
  assign __fsm_gemm_impl_in_state_15 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_15_index;
  assign __fsm_gemm_impl_in_state_7 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_7_index;
  assign __fsm_gemm_impl_in_state_14 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_14_index;
  assign __fsm_gemm_impl_in_state_6 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_6_index;
  assign and_11897 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_16;
  assign and_11898 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_8;
  assign __fsm_gemm_impl_in_state_12 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_12_index;
  assign __fsm_gemm_impl_in_state_4 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_4_index;
  assign ____fsm_gemm_impl_state__next_value_predicates = {nor_11679, __fsm_gemm_impl_returns_this_activation_vars};
  assign ____fsm___for_5_loop_state_0__next_value_predicates = {nor_11636, __fsm___for_5_loop_returns_this_activation_vars};
  assign p1_data_enable = p1_enable & p1_stage_done;
  assign p1_not_valid = ~p0_valid;
  assign p0_all_active_inputs_valid = (~__for_2_loop_contents_condition | v1_in_vld) & (~__for_1_loop_contents_condition | v0_in_vld);
  assign p0_all_active_outputs_ready = (~__for_2_loop_contents_condition | v1__write_req_rdy | __v1__write_req_has_been_sent_reg) & (v0__read_req_not_pred | v0__read_req_rdy | __v0__read_req_has_been_sent_reg) & (v0__read_req_not_pred | v1__read_req_rdy | __v1__read_req_has_been_sent_reg) & (~__for_1_loop_contents_condition | v0__write_req_rdy | __v0__write_req_has_been_sent_reg);
  assign __fsm_gemm_impl_in_state_2 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_2_index;
  assign __fsm_gemm_impl_in_state_3 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_3_index;
  assign __fsm_gemm_impl_in_state_5 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_5_index;
  assign __fsm_gemm_impl_in_state_9 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_9_index;
  assign __fsm_gemm_impl_in_state_10 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_10_index;
  assign __fsm_gemm_impl_in_state_11 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_11_index;
  assign __fsm_gemm_impl_in_state_13 = p1_____fsm_gemm_impl_state__1 == __fsm_gemm_impl_state_13_index;
  assign and_11905 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_15;
  assign and_11906 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_7;
  assign and_11907 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_14;
  assign and_11908 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_6;
  assign or_11910 = and_11897 | and_11898;
  assign and_11911 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_12;
  assign and_11912 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_4;
  assign C_ram_zero_latency0_select = __C_ram_zero_latency0_valid_skid_reg ? __C_ram_zero_latency0_skid_reg : C_rd_data;
  assign one_hot_11692 = {____fsm_gemm_impl_state__next_value_predicates[1:0] == 2'h0, ____fsm_gemm_impl_state__next_value_predicates[1] && !____fsm_gemm_impl_state__next_value_predicates[0], ____fsm_gemm_impl_state__next_value_predicates[0]};
  assign one_hot_11693 = {____fsm___for_5_loop_state_0__next_value_predicates[1:0] == 2'h0, ____fsm___for_5_loop_state_0__next_value_predicates[1] && !____fsm___for_5_loop_state_0__next_value_predicates[0], ____fsm___for_5_loop_state_0__next_value_predicates[0]};
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign p0_stage_done = p0_all_active_inputs_valid & p0_all_active_outputs_ready;
  assign and_11953 = p1_ctx_5__full_condition_ctx_6__ful_output & p1___fsm_gemm_impl_in_state_1;
  assign and_11924 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_2;
  assign and_11923 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_3;
  assign and_11921 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_5;
  assign and_11918 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_9;
  assign and_11917 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_10;
  assign and_11916 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_11;
  assign and_11915 = p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_13;
  assign or_11919 = and_11905 | and_11906;
  assign or_11920 = and_11907 | and_11908;
  assign or_11922 = or_11910 | and_11911 | and_11912;
  assign concat_11626 = {__fsm___for_5_loop_default_next_state, and_11582[2]};
  assign p0_data_enable = p0_enable & p0_stage_done;
  assign __v1__write_req_vld_buf = p0_all_active_inputs_valid & p0_enable & __for_2_loop_contents_condition;
  assign __v1__write_req_not_has_been_sent = ~__v1__write_req_has_been_sent_reg;
  assign __v0__read_req_vld_buf = p0_all_active_inputs_valid & p0_enable & nor_11636;
  assign __v0__read_req_not_has_been_sent = ~__v0__read_req_has_been_sent_reg;
  assign __v1__read_req_not_has_been_sent = ~__v1__read_req_has_been_sent_reg;
  assign __v0__write_req_vld_buf = p0_all_active_inputs_valid & p0_enable & __for_1_loop_contents_condition;
  assign __v0__write_req_not_has_been_sent = ~__v0__write_req_has_been_sent_reg;
  assign __C__read_req_vld_buf = p1_all_active_inputs_valid & p0_valid & p1_enable & or_11828;
  assign __C__read_req_not_has_been_sent = ~__C__read_req_has_been_sent_reg;
  assign or_11957 = p1___fsm___for_5_loop_returns_this_activation_vars | and_11953 | and_11924 | and_11923 | and_11912 | and_11921 | and_11908 | and_11906 | and_11898 | and_11918 | and_11917 | and_11916 | and_11911 | and_11915 | and_11907 | and_11905 | and_11897;
  assign __out_vld_buf = or_12447 & p1_valid & p1___for_6_loop_contents_condition;
  assign __out_not_has_been_sent = ~__out_has_been_sent_reg;
  assign and_12307 = p2_stage_done & p1_or_11828;
  assign C_write_value__16 = ____fsm___for_5_loop_state_3 + p1_smul_11826;
  assign C__read_resp_select = p1_or_11828 ? {C_ram_zero_latency0_select} : literal_11959;
  assign add_11673 = and_11590[1:0] + {__fsm___for_5_loop_default_next_state, and_11575[2]};
  assign add_11674 = and_11575[1:0] + concat_11626;
  assign __for_6_loop_contents_condition = __fsm_gemm_impl_in_state_18 & ctx_6__full_condition_continuati_output;
  assign add_11638 = and_11590[1:0] + concat_11626;
  assign and_12238 = nor_11679 & p0_data_enable;
  assign and_12239 = __fsm_gemm_impl_returns_this_activation_vars & p0_data_enable;
  assign and_12293 = nor_11636 & p0_data_enable;
  assign and_12294 = __fsm___for_5_loop_returns_this_activation_vars & p0_data_enable;
  assign __v1__write_req_valid_and_not_has_been_sent = __v1__write_req_vld_buf & __v1__write_req_not_has_been_sent;
  assign __v0__read_req_valid_and_not_has_been_sent = __v0__read_req_vld_buf & __v0__read_req_not_has_been_sent;
  assign __v1__read_req_valid_and_not_has_been_sent = __v0__read_req_vld_buf & __v1__read_req_not_has_been_sent;
  assign __v0__write_req_valid_and_not_has_been_sent = __v0__write_req_vld_buf & __v0__write_req_not_has_been_sent;
  assign C_rd_en__1 = __C__read_req_vld_buf & __C__read_req_not_has_been_sent;
  assign __C__write_req_vld_buf = or_12447 & p1_valid & or_11957;
  assign __C__write_req_not_has_been_sent = ~__C__write_req_has_been_sent_reg;
  assign __out_valid_and_not_has_been_sent = __out_vld_buf & __out_not_has_been_sent;
  assign C_ram_zero_latency0_to_is_not_rdy = ~and_12307;
  assign tuple_index_11964 = C__read_resp_select[31:0];
  assign v0_read_addr = {add_11673, and_11575[1:0]};
  assign v0_write_addr = and_11597[3:0];
  assign v0_in_select = __for_1_loop_contents_condition ? v0_in : 32'h0000_0000;
  assign v1_read_addr = {add_11674, and_11582[1:0]};
  assign v1_write_addr = and_11589[3:0];
  assign v1_in_select = __for_2_loop_contents_condition ? v1_in : 32'h0000_0000;
  assign ____fsm_gemm_impl_state__at_most_one_next_value = nor_11679 == one_hot_11692[1] & __fsm_gemm_impl_returns_this_activation_vars == one_hot_11692[0];
  assign ____fsm___for_5_loop_state_0__at_most_one_next_value = nor_11636 == one_hot_11693[1] & __fsm___for_5_loop_returns_this_activation_vars == one_hot_11693[0];
  assign concat_11648 = {nor_11636, __for_6_loop_contents_condition};
  assign C_read_addr__1 = and_11596[3:0];
  assign C_read_addr = {add_11638, and_11582[1:0]};
  assign concat_12241 = {and_12238, and_12239};
  assign __fsm_gemm_impl_state_plus_one = ____fsm_gemm_impl_state + __fsm_gemm_impl_state_1_index;
  assign v0__read_resp_select = p0_nor_11636 ? v0__read_resp : literal_11836;
  assign v1__read_resp_select = p0_nor_11636 ? v1__read_resp : literal_11840;
  assign continuation_1_ctx_3__full_condi_output = ~(__this[0] | __this[1]);
  assign __for_1_initial_loop_cond = ~and_11597[4];
  assign __for_2_guarded_update_state_elements = ~(~__fsm_gemm_impl_in_state_1 | ~ctx_5__full_condition_continuati_output | and_11589[4]);
  assign __for_3_initial_loop_cond = ~and_11590[2];
  assign __for_4_initial_loop_cond = ~and_11582[2];
  assign __for_5_initial_loop_cond = ~and_11575[2];
  assign __for_6_guarded_update_state_elements = ~(~__fsm_gemm_impl_in_state_18 | ~ctx_6__full_condition_continuati_output | and_11596[4]);
  assign concat_12296 = {and_12293, and_12294};
  assign __v1__write_req_valid_and_all_active_outputs_ready = __v1__write_req_vld_buf & p0_all_active_outputs_ready;
  assign __v1__write_req_valid_and_ready_txfr = __v1__write_req_valid_and_not_has_been_sent & v1__write_req_rdy;
  assign __v0__read_req_valid_and_all_active_outputs_ready = __v0__read_req_vld_buf & p0_all_active_outputs_ready;
  assign __v0__read_req_valid_and_ready_txfr = __v0__read_req_valid_and_not_has_been_sent & v0__read_req_rdy;
  assign __v1__read_req_valid_and_ready_txfr = __v1__read_req_valid_and_not_has_been_sent & v1__read_req_rdy;
  assign __v0__write_req_valid_and_all_active_outputs_ready = __v0__write_req_vld_buf & p0_all_active_outputs_ready;
  assign __v0__write_req_valid_and_ready_txfr = __v0__write_req_valid_and_not_has_been_sent & v0__write_req_rdy;
  assign __C__read_req_valid_and_all_active_outputs_ready = __C__read_req_vld_buf & or_12453;
  assign __C__read_req_valid_and_ready_txfr = C_rd_en__1 & C_ram_zero_latency0_from_skid_rdy;
  assign __C__write_req_valid_and_all_active_outputs_ready = __C__write_req_vld_buf & p2_all_active_outputs_ready;
  assign C_wr_en__1 = __C__write_req_vld_buf & __C__write_req_not_has_been_sent;
  assign __out_valid_and_all_active_outputs_ready = __out_vld_buf & p2_all_active_outputs_ready;
  assign __out_valid_and_ready_txfr = __out_valid_and_not_has_been_sent & out_rdy;
  assign C_ram_zero_latency0_skid_data_load_en = __C_rd_en__1_delay_reg & C_ram_zero_latency0_from_skid_rdy & C_ram_zero_latency0_to_is_not_rdy;
  assign C_ram_zero_latency0_skid_valid_set_zero = __C_ram_zero_latency0_valid_skid_reg & and_12307;
  assign tuple_11807 = {p0_tuple_11671_index0};
  assign tuple_11956 = {{and_11897 | and_11905 | and_11907 | and_11915 | and_11911 | and_11916 | and_11917 | and_11918 | p1_and_11664, or_11910 | or_11919 | or_11920 | and_11915 | and_11921 | p1_and_11665, or_11922 | or_11919 | and_11916 | and_11923 | p1_and_11666, or_11922 | or_11920 | and_11917 | and_11924 | p1_and_11667}, C_write_value__16 & {32{p1___fsm___for_5_loop_returns_this_activation_vars}}};
  assign C_read_response__1 = tuple_index_11964 & {32{p1___for_6_loop_contents_condition}};
  assign and_12309 = p1_data_enable & p0_nor_11636;
  assign and_12311 = p0_data_enable & __for_1_loop_contents_condition;
  assign and_12314 = p0_data_enable & __for_2_loop_contents_condition;
  assign or_12444 = ~p0_stage_done | ____fsm_gemm_impl_state__at_most_one_next_value | rst;
  assign or_12446 = ~p0_stage_done | ____fsm___for_5_loop_state_0__at_most_one_next_value | rst;
  assign p3_enable = 1'h1;
  assign p2_enable = 1'h1;
  assign nand_11970 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & p1___fsm_gemm_impl_in_state_1);
  assign nand_11971 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_2);
  assign nand_11972 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_3);
  assign nand_11973 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_4);
  assign nand_11974 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_5);
  assign nand_11975 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_6);
  assign nand_11976 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_7);
  assign nand_11977 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_8);
  assign nand_11978 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_9);
  assign nand_11979 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_10);
  assign nand_11980 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_11);
  assign nand_11981 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_12);
  assign nand_11982 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_13);
  assign nand_11983 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_14);
  assign nand_11984 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_15);
  assign nand_11985 = ~(p1_ctx_5__full_condition_ctx_6__ful_output & __fsm_gemm_impl_in_state_16);
  assign smul_11826 = smul32b_32b_x_32b(____fsm___for_5_loop_state_1, ____fsm___for_5_loop_state_2);
  assign one_hot_sel_11662 = C_read_addr__1 & {4{concat_11648[0]}} | C_read_addr & {4{concat_11648[1]}};
  assign nand_11745 = ~(~ne_11602 & ctx_5__full_condition_ctx_6__ful_output & ____fsm___for_5_loop_state_0);
  assign nand_11746 = ~(__fsm_gemm_impl_in_state_18 & ctx_6__full_condition_continuati_output);
  assign nand_11747 = ~(~ne_11602 & ctx_5__full_condition_ctx_6__ful_output & __fsm___for_5_loop_in_state_0);
  assign and_11664 = __fsm___for_5_loop_returns_this_activation_vars & add_11638[1];
  assign and_11665 = __fsm___for_5_loop_returns_this_activation_vars & add_11638[0];
  assign and_11666 = __fsm___for_5_loop_returns_this_activation_vars & and_11582[1];
  assign and_11667 = __fsm___for_5_loop_returns_this_activation_vars & and_11582[0];
  assign one_hot_sel_12242 = __fsm_gemm_impl_state_0_index & {5{concat_12241[0]}} | __fsm_gemm_impl_state_plus_one & {5{concat_12241[1]}};
  assign or_12243 = and_12238 | and_12239;
  assign and_12251 = __for_4_do_break_with_fsm & p0_data_enable;
  assign and_12254 = __for_5_do_break_with_fsm & p0_data_enable;
  assign v0_read_response = v0__read_resp_select[31:0];
  assign and_12260 = p0___fsm___for_5_loop_in_state_0 & p1_data_enable;
  assign v1_read_response = v1__read_resp_select[31:0];
  assign C_read_response = tuple_index_11964 & {32{p1_nor_11636}};
  assign and_12266 = p1___fsm___for_5_loop_in_state_0 & p2_stage_done;
  assign and_12269 = __for_6_loop_contents_condition & p0_data_enable;
  assign unexpand_for_this_next__1_case_1 = literal_11493[__this];
  assign unexpand_for___for_1__i_next__1_case_1 = add_11617[4:0];
  assign and_12463 = __fsm_gemm_impl_in_state_0 & continuation_1_ctx_3__full_condi_output & __for_1_initial_loop_cond & p0_data_enable;
  assign unexpand_for___for_2__i_next__1_case_1 = add_11609[4:0];
  assign and_12278 = __for_2_guarded_update_state_elements & p0_data_enable;
  assign unexpand_for___for_3_i_next__1_case_1 = add_11610[2:0];
  assign and_12464 = __for_4_do_break_with_fsm & __for_3_initial_loop_cond & p0_data_enable;
  assign unexpand_for___for_4_j_next__1_case_1 = add_11600[2:0];
  assign and_12465 = __for_5_do_break_with_fsm & __for_4_initial_loop_cond & p0_data_enable;
  assign unexpand_for___for_5_k_next__1_case_1 = add_11592[2:0];
  assign and_12466 = __fsm___for_5_loop_returns_this_activation_vars & __for_5_initial_loop_cond & p0_data_enable;
  assign unexpand_for___for_6__i_next__1_case_1 = add_11614[4:0];
  assign and_12290 = __for_6_guarded_update_state_elements & p0_data_enable;
  assign one_hot_sel_12297 = __fsm___for_5_loop_default_next_state & concat_12296[0] | __for_4_enter_condition & concat_12296[1];
  assign or_12298 = and_12293 | and_12294;
  assign __v1__write_req_not_stage_load = ~__v1__write_req_valid_and_all_active_outputs_ready;
  assign __v1__write_req_has_been_sent_reg_load_en = __v1__write_req_valid_and_ready_txfr | __v1__write_req_valid_and_all_active_outputs_ready;
  assign __v0__read_req_not_stage_load = ~__v0__read_req_valid_and_all_active_outputs_ready;
  assign __v0__read_req_has_been_sent_reg_load_en = __v0__read_req_valid_and_ready_txfr | __v0__read_req_valid_and_all_active_outputs_ready;
  assign __v1__read_req_has_been_sent_reg_load_en = __v1__read_req_valid_and_ready_txfr | __v0__read_req_valid_and_all_active_outputs_ready;
  assign __v0__write_req_not_stage_load = ~__v0__write_req_valid_and_all_active_outputs_ready;
  assign __v0__write_req_has_been_sent_reg_load_en = __v0__write_req_valid_and_ready_txfr | __v0__write_req_valid_and_all_active_outputs_ready;
  assign __C__read_req_not_stage_load = ~__C__read_req_valid_and_all_active_outputs_ready;
  assign __C__read_req_has_been_sent_reg_load_en = __C__read_req_valid_and_ready_txfr | __C__read_req_valid_and_all_active_outputs_ready;
  assign __C__write_req_not_stage_load = ~__C__write_req_valid_and_all_active_outputs_ready;
  assign __C__write_req_has_been_sent_reg_load_en = C_wr_en__1 | __C__write_req_valid_and_all_active_outputs_ready;
  assign __out_not_stage_load = ~__out_valid_and_all_active_outputs_ready;
  assign __out_has_been_sent_reg_load_en = __out_valid_and_ready_txfr | __out_valid_and_all_active_outputs_ready;
  assign C_ram_zero_latency0_skid_valid_load_en = C_ram_zero_latency0_skid_data_load_en | C_ram_zero_latency0_skid_valid_set_zero;
  always_ff @ (posedge clk) begin
    if (rst) begin
      ____for_5__last_iter_broke <= 1'h1;
      ____for_4__last_iter_broke <= 1'h1;
      ____for_2__last_iter_broke <= 1'h1;
      ____for_3__last_iter_broke <= 1'h1;
      ____for_5_k <= 3'h0;
      ____for_6__last_iter_broke <= 1'h1;
      ____for_1__last_iter_broke <= 1'h1;
      ____for_4_j <= 3'h0;
      ____for_2__i <= 5'h00;
      ____for_3_i <= 3'h0;
      __this <= 2'h0;
      ____for_6__i <= 5'h00;
      ____for_1__i <= 5'h00;
      ____fsm_gemm_impl_state <= 5'h00;
      ____fsm___for_5_loop_state_0 <= 1'h0;
      p0_____fsm_gemm_impl_state__1 <= 5'h00;
      p0_____fsm___for_5_loop_state_0__1 <= 1'h0;
      p0___fsm_gemm_impl_in_state_1 <= 1'h0;
      p0___for_2_loop_contents_condition <= 1'h0;
      p0_ctx_5__full_condition_ctx_6__ful_output <= 1'h0;
      p0___fsm___for_5_loop_in_state_0 <= 1'h0;
      p0___fsm___for_5_loop_returns_this_activation_vars <= 1'h0;
      p0___for_6_loop_contents_condition <= 1'h0;
      p0_nor_11636 <= 1'h0;
      p0___for_1_loop_contents_condition <= 1'h0;
      p0_tuple_11671_index0 <= 4'h0;
      p0_nand_11745 <= 1'h0;
      p0_nand_11746 <= 1'h0;
      p0_nand_11747 <= 1'h0;
      p0_and_11664 <= 1'h0;
      p0_and_11665 <= 1'h0;
      p0_and_11666 <= 1'h0;
      p0_and_11667 <= 1'h0;
      ____fsm___for_5_loop_state_1 <= 32'h0000_0000;
      ____fsm___for_5_loop_state_2 <= 32'h0000_0000;
      p1_____fsm_gemm_impl_state__1 <= 5'h00;
      p1_____fsm___for_5_loop_state_0__1 <= 1'h0;
      p1___fsm_gemm_impl_in_state_1 <= 1'h0;
      p1_ctx_5__full_condition_ctx_6__ful_output <= 1'h0;
      p1___fsm___for_5_loop_in_state_0 <= 1'h0;
      p1___fsm___for_5_loop_returns_this_activation_vars <= 1'h0;
      p1_smul_11826 <= 32'h0000_0000;
      p1___for_6_loop_contents_condition <= 1'h0;
      p1_nor_11636 <= 1'h0;
      p1_or_11828 <= 1'h0;
      p1_nand_11745 <= 1'h0;
      p1_nand_11746 <= 1'h0;
      p1_nand_11747 <= 1'h0;
      p1_and_11664 <= 1'h0;
      p1_and_11665 <= 1'h0;
      p1_and_11666 <= 1'h0;
      p1_and_11667 <= 1'h0;
      ____fsm___for_5_loop_state_3 <= 32'h0000_0000;
      p2___fsm___for_5_loop_returns_this_activation_vars <= 1'h0;
      p2_and_11953 <= 1'h0;
      p2_and_11924 <= 1'h0;
      p2_and_11923 <= 1'h0;
      p2_and_11912 <= 1'h0;
      p2_and_11921 <= 1'h0;
      p2_and_11908 <= 1'h0;
      p2_and_11906 <= 1'h0;
      p2_and_11898 <= 1'h0;
      p2_and_11918 <= 1'h0;
      p2_and_11917 <= 1'h0;
      p2_and_11916 <= 1'h0;
      p2_and_11911 <= 1'h0;
      p2_and_11915 <= 1'h0;
      p2_and_11907 <= 1'h0;
      p2_and_11905 <= 1'h0;
      p2_and_11897 <= 1'h0;
      p2_or_11957 <= 1'h0;
      p2_nand_11745 <= 1'h0;
      p2_nand_11970 <= 1'h0;
      p2_nand_11971 <= 1'h0;
      p2_nand_11972 <= 1'h0;
      p2_nand_11973 <= 1'h0;
      p2_nand_11974 <= 1'h0;
      p2_nand_11975 <= 1'h0;
      p2_nand_11976 <= 1'h0;
      p2_nand_11977 <= 1'h0;
      p2_nand_11978 <= 1'h0;
      p2_nand_11979 <= 1'h0;
      p2_nand_11980 <= 1'h0;
      p2_nand_11981 <= 1'h0;
      p2_nand_11982 <= 1'h0;
      p2_nand_11983 <= 1'h0;
      p2_nand_11984 <= 1'h0;
      p2_nand_11985 <= 1'h0;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      __v1__write_req_has_been_sent_reg <= 1'h0;
      __v0__read_req_has_been_sent_reg <= 1'h0;
      __v1__read_req_has_been_sent_reg <= 1'h0;
      __v0__write_req_has_been_sent_reg <= 1'h0;
      __C__read_req_has_been_sent_reg <= 1'h0;
      __C__write_req_has_been_sent_reg <= 1'h0;
      __out_has_been_sent_reg <= 1'h0;
      __C_rd_en__1_delay_reg <= 1'h0;
      __C_ram_zero_latency0_skid_reg <= 32'h0000_0000;
      __C_ram_zero_latency0_valid_skid_reg <= 1'h0;
    end else begin
      ____for_5__last_iter_broke <= and_12294 ? __for_5_do_break_from_func : ____for_5__last_iter_broke;
      ____for_4__last_iter_broke <= and_12254 ? __for_4_do_break_from_func : ____for_4__last_iter_broke;
      ____for_2__last_iter_broke <= and_12314 ? __for_2_do_break_from_func : ____for_2__last_iter_broke;
      ____for_3__last_iter_broke <= and_12251 ? __for_3_do_break_from_func : ____for_3__last_iter_broke;
      ____for_5_k <= and_12466 ? unexpand_for___for_5_k_next__1_case_1 : ____for_5_k;
      ____for_6__last_iter_broke <= and_12269 ? __for_6_do_break_from_func : ____for_6__last_iter_broke;
      ____for_1__last_iter_broke <= and_12311 ? __for_1_do_break_from_func : ____for_1__last_iter_broke;
      ____for_4_j <= and_12465 ? unexpand_for___for_4_j_next__1_case_1 : ____for_4_j;
      ____for_2__i <= and_12278 ? unexpand_for___for_2__i_next__1_case_1 : ____for_2__i;
      ____for_3_i <= and_12464 ? unexpand_for___for_3_i_next__1_case_1 : ____for_3_i;
      __this <= and_12239 ? unexpand_for_this_next__1_case_1 : __this;
      ____for_6__i <= and_12290 ? unexpand_for___for_6__i_next__1_case_1 : ____for_6__i;
      ____for_1__i <= and_12463 ? unexpand_for___for_1__i_next__1_case_1 : ____for_1__i;
      ____fsm_gemm_impl_state <= or_12243 ? one_hot_sel_12242 : ____fsm_gemm_impl_state;
      ____fsm___for_5_loop_state_0 <= or_12298 ? one_hot_sel_12297 : ____fsm___for_5_loop_state_0;
      p0_____fsm_gemm_impl_state__1 <= p0_data_enable ? ____fsm_gemm_impl_state : p0_____fsm_gemm_impl_state__1;
      p0_____fsm___for_5_loop_state_0__1 <= p0_data_enable ? ____fsm___for_5_loop_state_0 : p0_____fsm___for_5_loop_state_0__1;
      p0___fsm_gemm_impl_in_state_1 <= p0_data_enable ? __fsm_gemm_impl_in_state_1 : p0___fsm_gemm_impl_in_state_1;
      p0___for_2_loop_contents_condition <= p0_data_enable ? __for_2_loop_contents_condition : p0___for_2_loop_contents_condition;
      p0_ctx_5__full_condition_ctx_6__ful_output <= p0_data_enable ? ctx_5__full_condition_ctx_6__ful_output : p0_ctx_5__full_condition_ctx_6__ful_output;
      p0___fsm___for_5_loop_in_state_0 <= p0_data_enable ? __fsm___for_5_loop_in_state_0 : p0___fsm___for_5_loop_in_state_0;
      p0___fsm___for_5_loop_returns_this_activation_vars <= p0_data_enable ? __fsm___for_5_loop_returns_this_activation_vars : p0___fsm___for_5_loop_returns_this_activation_vars;
      p0___for_6_loop_contents_condition <= p0_data_enable ? __for_6_loop_contents_condition : p0___for_6_loop_contents_condition;
      p0_nor_11636 <= p0_data_enable ? nor_11636 : p0_nor_11636;
      p0___for_1_loop_contents_condition <= p0_data_enable ? __for_1_loop_contents_condition : p0___for_1_loop_contents_condition;
      p0_tuple_11671_index0 <= p0_data_enable ? one_hot_sel_11662 : p0_tuple_11671_index0;
      p0_nand_11745 <= p0_data_enable ? nand_11745 : p0_nand_11745;
      p0_nand_11746 <= p0_data_enable ? nand_11746 : p0_nand_11746;
      p0_nand_11747 <= p0_data_enable ? nand_11747 : p0_nand_11747;
      p0_and_11664 <= p0_data_enable ? and_11664 : p0_and_11664;
      p0_and_11665 <= p0_data_enable ? and_11665 : p0_and_11665;
      p0_and_11666 <= p0_data_enable ? and_11666 : p0_and_11666;
      p0_and_11667 <= p0_data_enable ? and_11667 : p0_and_11667;
      ____fsm___for_5_loop_state_1 <= and_12260 ? v0_read_response : ____fsm___for_5_loop_state_1;
      ____fsm___for_5_loop_state_2 <= and_12260 ? v1_read_response : ____fsm___for_5_loop_state_2;
      p1_____fsm_gemm_impl_state__1 <= p1_data_enable ? p0_____fsm_gemm_impl_state__1 : p1_____fsm_gemm_impl_state__1;
      p1_____fsm___for_5_loop_state_0__1 <= p1_data_enable ? p0_____fsm___for_5_loop_state_0__1 : p1_____fsm___for_5_loop_state_0__1;
      p1___fsm_gemm_impl_in_state_1 <= p1_data_enable ? p0___fsm_gemm_impl_in_state_1 : p1___fsm_gemm_impl_in_state_1;
      p1_ctx_5__full_condition_ctx_6__ful_output <= p1_data_enable ? p0_ctx_5__full_condition_ctx_6__ful_output : p1_ctx_5__full_condition_ctx_6__ful_output;
      p1___fsm___for_5_loop_in_state_0 <= p1_data_enable ? p0___fsm___for_5_loop_in_state_0 : p1___fsm___for_5_loop_in_state_0;
      p1___fsm___for_5_loop_returns_this_activation_vars <= p1_data_enable ? p0___fsm___for_5_loop_returns_this_activation_vars : p1___fsm___for_5_loop_returns_this_activation_vars;
      p1_smul_11826 <= p1_data_enable ? smul_11826 : p1_smul_11826;
      p1___for_6_loop_contents_condition <= p1_data_enable ? p0___for_6_loop_contents_condition : p1___for_6_loop_contents_condition;
      p1_nor_11636 <= p1_data_enable ? p0_nor_11636 : p1_nor_11636;
      p1_or_11828 <= p1_data_enable ? or_11828 : p1_or_11828;
      p1_nand_11745 <= p1_data_enable ? p0_nand_11745 : p1_nand_11745;
      p1_nand_11746 <= p1_data_enable ? p0_nand_11746 : p1_nand_11746;
      p1_nand_11747 <= p1_data_enable ? p0_nand_11747 : p1_nand_11747;
      p1_and_11664 <= p1_data_enable ? p0_and_11664 : p1_and_11664;
      p1_and_11665 <= p1_data_enable ? p0_and_11665 : p1_and_11665;
      p1_and_11666 <= p1_data_enable ? p0_and_11666 : p1_and_11666;
      p1_and_11667 <= p1_data_enable ? p0_and_11667 : p1_and_11667;
      ____fsm___for_5_loop_state_3 <= and_12266 ? C_read_response : ____fsm___for_5_loop_state_3;
      p2___fsm___for_5_loop_returns_this_activation_vars <= p2_stage_done ? p1___fsm___for_5_loop_returns_this_activation_vars : p2___fsm___for_5_loop_returns_this_activation_vars;
      p2_and_11953 <= p2_stage_done ? and_11953 : p2_and_11953;
      p2_and_11924 <= p2_stage_done ? and_11924 : p2_and_11924;
      p2_and_11923 <= p2_stage_done ? and_11923 : p2_and_11923;
      p2_and_11912 <= p2_stage_done ? and_11912 : p2_and_11912;
      p2_and_11921 <= p2_stage_done ? and_11921 : p2_and_11921;
      p2_and_11908 <= p2_stage_done ? and_11908 : p2_and_11908;
      p2_and_11906 <= p2_stage_done ? and_11906 : p2_and_11906;
      p2_and_11898 <= p2_stage_done ? and_11898 : p2_and_11898;
      p2_and_11918 <= p2_stage_done ? and_11918 : p2_and_11918;
      p2_and_11917 <= p2_stage_done ? and_11917 : p2_and_11917;
      p2_and_11916 <= p2_stage_done ? and_11916 : p2_and_11916;
      p2_and_11911 <= p2_stage_done ? and_11911 : p2_and_11911;
      p2_and_11915 <= p2_stage_done ? and_11915 : p2_and_11915;
      p2_and_11907 <= p2_stage_done ? and_11907 : p2_and_11907;
      p2_and_11905 <= p2_stage_done ? and_11905 : p2_and_11905;
      p2_and_11897 <= p2_stage_done ? and_11897 : p2_and_11897;
      p2_or_11957 <= p2_stage_done ? or_11957 : p2_or_11957;
      p2_nand_11745 <= p2_stage_done ? p1_nand_11745 : p2_nand_11745;
      p2_nand_11970 <= p2_stage_done ? nand_11970 : p2_nand_11970;
      p2_nand_11971 <= p2_stage_done ? nand_11971 : p2_nand_11971;
      p2_nand_11972 <= p2_stage_done ? nand_11972 : p2_nand_11972;
      p2_nand_11973 <= p2_stage_done ? nand_11973 : p2_nand_11973;
      p2_nand_11974 <= p2_stage_done ? nand_11974 : p2_nand_11974;
      p2_nand_11975 <= p2_stage_done ? nand_11975 : p2_nand_11975;
      p2_nand_11976 <= p2_stage_done ? nand_11976 : p2_nand_11976;
      p2_nand_11977 <= p2_stage_done ? nand_11977 : p2_nand_11977;
      p2_nand_11978 <= p2_stage_done ? nand_11978 : p2_nand_11978;
      p2_nand_11979 <= p2_stage_done ? nand_11979 : p2_nand_11979;
      p2_nand_11980 <= p2_stage_done ? nand_11980 : p2_nand_11980;
      p2_nand_11981 <= p2_stage_done ? nand_11981 : p2_nand_11981;
      p2_nand_11982 <= p2_stage_done ? nand_11982 : p2_nand_11982;
      p2_nand_11983 <= p2_stage_done ? nand_11983 : p2_nand_11983;
      p2_nand_11984 <= p2_stage_done ? nand_11984 : p2_nand_11984;
      p2_nand_11985 <= p2_stage_done ? nand_11985 : p2_nand_11985;
      p0_valid <= p0_enable ? p0_stage_done : p0_valid;
      p1_valid <= p1_enable ? p1_stage_done : p1_valid;
      p2_valid <= p2_enable ? p2_stage_done : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      __v1__write_req_has_been_sent_reg <= __v1__write_req_has_been_sent_reg_load_en ? __v1__write_req_not_stage_load : __v1__write_req_has_been_sent_reg;
      __v0__read_req_has_been_sent_reg <= __v0__read_req_has_been_sent_reg_load_en ? __v0__read_req_not_stage_load : __v0__read_req_has_been_sent_reg;
      __v1__read_req_has_been_sent_reg <= __v1__read_req_has_been_sent_reg_load_en ? __v0__read_req_not_stage_load : __v1__read_req_has_been_sent_reg;
      __v0__write_req_has_been_sent_reg <= __v0__write_req_has_been_sent_reg_load_en ? __v0__write_req_not_stage_load : __v0__write_req_has_been_sent_reg;
      __C__read_req_has_been_sent_reg <= __C__read_req_has_been_sent_reg_load_en ? __C__read_req_not_stage_load : __C__read_req_has_been_sent_reg;
      __C__write_req_has_been_sent_reg <= __C__write_req_has_been_sent_reg_load_en ? __C__write_req_not_stage_load : __C__write_req_has_been_sent_reg;
      __out_has_been_sent_reg <= __out_has_been_sent_reg_load_en ? __out_not_stage_load : __out_has_been_sent_reg;
      __C_rd_en__1_delay_reg <= C_rd_en__1;
      __C_ram_zero_latency0_skid_reg <= C_ram_zero_latency0_skid_data_load_en ? C_rd_data : __C_ram_zero_latency0_skid_reg;
      __C_ram_zero_latency0_valid_skid_reg <= C_ram_zero_latency0_skid_valid_load_en ? C_ram_zero_latency0_from_skid_rdy : __C_ram_zero_latency0_valid_skid_reg;
    end
  end
  assign out = C_read_response__1;
  assign out_vld = __out_valid_and_not_has_been_sent;
  assign v0__read_req = {v0_read_addr};
  assign v0__read_req_vld = __v0__read_req_valid_and_not_has_been_sent;
  assign v0__read_resp_rdy = and_12309;
  assign v0__write_completion_rdy = p1_data_enable & p0___for_1_loop_contents_condition;
  assign v0__write_req = {v0_write_addr, v0_in_select};
  assign v0__write_req_vld = __v0__write_req_valid_and_not_has_been_sent;
  assign v0_in_rdy = and_12311;
  assign v1__read_req = {v1_read_addr};
  assign v1__read_req_vld = __v1__read_req_valid_and_not_has_been_sent;
  assign v1__read_resp_rdy = and_12309;
  assign v1__write_completion_rdy = p1_data_enable & p0___for_2_loop_contents_condition;
  assign v1__write_req = {v1_write_addr, v1_in_select};
  assign v1__write_req_vld = __v1__write_req_valid_and_not_has_been_sent;
  assign v1_in_rdy = and_12314;
  assign C_rd_addr = tuple_11807[3:0];
  assign C_rd_en = C_rd_en__1;
  assign C_wr_addr = tuple_11956[35:32];
  assign C_wr_data = tuple_11956[31:0];
  assign C_wr_en = C_wr_en__1;
  `ifdef ASSERT_ON
  ____fsm_gemm_impl_state__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_12444))) or_12444) else $fatal(0, "More than one next_value fired for state element: __fsm_gemm_impl_state");
  ____fsm___for_5_loop_state_0__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_12446))) or_12446) else $fatal(0, "More than one next_value fired for state element: __fsm___for_5_loop_state_0");
  `endif  // ASSERT_ON
endmodule
